module ACC54(SFTCTRL, DSPIN, PP, CINPUT, LOAD, M9ADDSUB, ADDSUB, CIN, CASIN, CEO, RSTO, CEC, RSTC, CLK, SIGNEDI, SUM1, SUM0, DSPOUT, CASCOUT, ROUNDEN, CECIN, CECTRL, RSTCIN, RSTCTRL); //synthesis syn_black_box syn_lib_cell=1
    input [3:0] SFTCTRL;
    input [53:0] DSPIN;
    input [71:0] PP;
    input [53:0] CINPUT;
    input LOAD;
    input [1:0] M9ADDSUB;
    input [1:0] ADDSUB;
    input CIN;
    input [1:0] CASIN;
    input CEO;
    input RSTO;
    input CEC;
    input RSTC;
    input CLK;
    input SIGNEDI;
    output [35:0] SUM1;
    output [35:0] SUM0;
    output [53:0] DSPOUT;
    output [1:0] CASCOUT;
    input ROUNDEN;
    input CECIN;
    input CECTRL;
    input RSTCIN;
    input RSTCTRL;
    parameter SIGN = "DISABLED";
    parameter M9ADDSUB_CTRL = "ADDITION";
    parameter ADDSUB_CTRL = "ADD_ADD_CTRL_54_BIT_ADDER";
    parameter STATICOPCODE_EN = "DISABLED";
    parameter OUTREGBYPS = "REGISTER";
    parameter GSR = "ENABLED";
    parameter PROGCONST = "0b000000000000000000000000000000000000000000000000000000";
    parameter CONSTSEL = "BYPASS";
    parameter DSPCASCADE = "DISABLED";
    parameter ACC108CASCADE = "BYPASSCASCADE";
    parameter ACCUMODE = "MODE0";
    parameter ACCUBYPS = "USED";
    parameter CREGBYPS1 = "REGISTER";
    parameter CREGBYPS2 = "REGISTER";
    parameter CREGBYPS3 = "REGISTER";
    parameter CINREGBYPS1 = "REGISTER";
    parameter CINREGBYPS2 = "REGISTER";
    parameter CINREGBYPS3 = "REGISTER";
    parameter LOADREGBYPS1 = "REGISTER";
    parameter LOADREGBYPS2 = "REGISTER";
    parameter LOADREGBYPS3 = "REGISTER";
    parameter M9ADDSUBREGBYPS1 = "REGISTER";
    parameter M9ADDSUBREGBYPS2 = "REGISTER";
    parameter M9ADDSUBREGBYPS3 = "REGISTER";
    parameter ADDSUBSIGNREGBYPS1 = "REGISTER";
    parameter ADDSUBSIGNREGBYPS2 = "REGISTER";
    parameter ADDSUBSIGNREGBYPS3 = "REGISTER";
    parameter ROUNDHALFUP = "DISABLED";
    parameter ROUNDRTZI = "ROUND_TO_ZERO";
    parameter ROUNDBIT = "ROUND_TO_BIT0";
    parameter CASCOUTREGBYPS = "REGISTER";
    parameter SFTEN = "DISABLED";
    parameter RESET = "SYNC";
endmodule

module ADC(DN0, DN1, DP0, DP1, ADCEN, CAL, CALRDY, CHAEN, CHASEL, CHBEN, CHBSEL, CLKDCLK, CLKFAB, COG, COMP1IN, COMP1IP, COMP1OL, COMP2IN, COMP2IP, COMP2OL, COMP3IN, COMP3IP, COMP3OL, CONVSTOP, DA, DB, EOC, GPION, GPIOP, RESETN, RSTN, SOC, COMP1O, COMP2O, COMP3O); //synthesis black_box_pad_pin="DN0,DN1,DP0,DP1" syn_lib_cell=1
    input DN0;
    input DN1;
    input DP0;
    input DP1;
    input ADCEN;
    input CAL;
    output CALRDY;
    input CHAEN;
    input [3:0] CHASEL;
    input CHBEN;
    input [3:0] CHBSEL;
    input CLKDCLK;
    input CLKFAB;
    output COG;
    input COMP1IN;
    input COMP1IP;
    output COMP1OL;
    input COMP2IN;
    input COMP2IP;
    output COMP2OL;
    input COMP3IN;
    input COMP3IP;
    output COMP3OL;
    input CONVSTOP;
    output [11:0] DA;
    output [11:0] DB;
    output EOC;
    input [15:0] GPION;
    input [15:0] GPIOP;
    input RESETN;
    input RSTN;
    input SOC;
    output COMP1O;
    output COMP2O;
    output COMP3O;
    parameter ADC_ENP = "ENABLED";
    parameter CLK_DIV = "2";
    parameter CTLCOMPSW1 = "DISABLED";
    parameter CTLCOMPSW2 = "DISABLED";
    parameter CTLCOMPSW3 = "DISABLED";
    parameter DF = "STRAIGHT_BINARY";
    parameter EN_COMP1 = "ENABLED";
    parameter EN_COMP2 = "ENABLED";
    parameter EN_COMP3 = "ENABLED";
    parameter OMA = "BIPOLAR";
    parameter OMB = "BIPOLAR";
    parameter REFBUFAEN = "ENABLED";
    parameter REFBUFBEN = "ENABLED";
    parameter SLEEP = "DISABLED";
    parameter VREFACFG = "1P0_TO_1P2";
    parameter VREFASEL = "INTERNAL";
    parameter VREFBCFG = "1P0_TO_1P2";
    parameter VREFBSEL = "INTERNAL";
endmodule

module ALUREG(ALUCLK, ALUFLAGC, ALUFLAGV, ALUFLAGZ, ALUFORWARDA, ALUFORWARDB, ALUIREGEN, ALUOREGEN, ALURST, DATAA, DATAB, DATAC, OPC, OPCCUSTOM, RADDRA, RADDRB, RDATAA, RDATAB, REGCLK, REGCLKEN, REGRST, RESULT, WADDR, WDROTATE, WDSIGNEXT, WDSIZE, WDATA, WREN); //synthesis syn_black_box syn_lib_cell=1
    input ALUCLK;
    output ALUFLAGC;
    output ALUFLAGV;
    output ALUFLAGZ;
    input ALUFORWARDA;
    input ALUFORWARDB;
    input ALUIREGEN;
    input ALUOREGEN;
    input ALURST;
    input [31:0] DATAA;
    input [31:0] DATAB;
    input [4:0] DATAC;
    input [6:0] OPC;
    input OPCCUSTOM;
    input [4:0] RADDRA;
    input [4:0] RADDRB;
    output [31:0] RDATAA;
    output [31:0] RDATAB;
    input REGCLK;
    input REGCLKEN;
    input REGRST;
    output [31:0] RESULT;
    input [4:0] WADDR;
    input [1:0] WDROTATE;
    input WDSIGNEXT;
    input [1:0] WDSIZE;
    input [31:0] WDATA;
    input WREN;
    parameter ALURST_ACTIVELOW = "DISABLE";
    parameter GSR = "ENABLED";
    parameter INREG = "DISABLE";
    parameter MULFXP_ROUND = "ENABLE";
    parameter OUTREG = "DISABLE";
    parameter REGRST_ACTIVELOW = "DISABLE";
    parameter RETAIN = "ENABLE";
    parameter RFASYNC_RD = "SYNC_RD";
    parameter RFR0_RO = "R0READONLY";
    parameter RFUNALIA_WR = "DISABLE";
    parameter RFWCLK_INV = "SIG";
endmodule

module BB_ADC(IOPAD, INADC); //synthesis black_box_pad_pin="IOPAD" syn_lib_cell=1
    inout IOPAD;
    output INADC;
endmodule

module BB_CDR(IOPAD, INADC); //synthesis black_box_pad_pin="IOPAD" syn_lib_cell=1
    inout IOPAD;
    output INADC;
endmodule

module BB_I3C_A(IOPAD, PADDI, PADDO, PADDT, I3CRESEN, I3CWKPU); //synthesis black_box_pad_pin="IOPAD" syn_lib_cell=1
    inout IOPAD;
    output PADDI;
    input PADDO;
    input PADDT;
    input I3CRESEN;
    input I3CWKPU;
endmodule

module BFD1P3KX(DOUT, DIN, DT, CEOUT, CLKOUT, SROUT, CEIN, CLKIN, SRIN, QOUT, QIN, QT); //synthesis syn_black_box syn_lib_cell=1
    input DOUT;
    input DIN;
    input DT;
    input CEOUT;
    input CLKOUT;
    input SROUT;
    input CEIN;
    input CLKIN;
    input SRIN;
    output QOUT;
    output QIN;
    output QT;
    parameter GSR = "ENABLED";
    parameter OUTSET = "RESET";
    parameter INSET = "RESET";
    parameter TSSET = "RESET";
endmodule

module BFD1P3LX(DOUT, DIN, DT, CEOUT, CLKOUT, SROUT, CEIN, CLKIN, SRIN, QOUT, QIN, QT); //synthesis syn_black_box syn_lib_cell=1
    input DOUT;
    input DIN;
    input DT;
    input CEOUT;
    input CLKOUT;
    input SROUT;
    input CEIN;
    input CLKIN;
    input SRIN;
    output QOUT;
    output QIN;
    output QT;
    parameter GSR = "ENABLED";
    parameter OUTSET = "RESET";
    parameter INSET = "RESET";
    parameter TSSET = "RESET";
endmodule

module BNKREF18(STDBYINR, STDBYDIF, PVTCODE); //synthesis syn_noprune=1 syn_lib_cell=1
    input STDBYINR;
    input STDBYDIF;
    output [6:0] PVTCODE;
    parameter BANK = "0b0000";
    parameter STANDBY_DIFFIO = "DISABLED";
    parameter STANDBY_INR = "DISABLED";
endmodule

module CONFIG_LMMI(LMMICLK, LMMIREQUEST, LMMIWRRD_N, LMMIOFFSET, LMMIWDATA, LMMIRDATA, LMMIREADY, LMMIRDATAVALID, LMMIRESETN, RSTSMCLK, SMCLK); //synthesis syn_black_box syn_lib_cell=1
    input LMMICLK;
    input LMMIREQUEST;
    input LMMIWRRD_N;
    input [7:0] LMMIOFFSET;
    input [7:0] LMMIWDATA;
    output [7:0] LMMIRDATA;
    output LMMIREADY;
    output LMMIRDATAVALID;
    input LMMIRESETN;
    input RSTSMCLK;
    input SMCLK;
    parameter LMMI_EN = "DIS";
endmodule

module DDRDLL(CODE, FREEZE, LOCK, CLKIN, RST, DCNTL, UDDCNTL_N); //synthesis syn_black_box syn_lib_cell=1
    output [8:0] CODE;
    input FREEZE;
    output LOCK;
    input CLKIN;
    input RST;
    output [8:0] DCNTL;
    input UDDCNTL_N;
    parameter GSR = "ENABLED";
    parameter ENA_ROUNDOFF = "ENABLED";
    parameter FORCE_MAX_DELAY = "CODE_OR_LOCK_FROM_DLL_LOOP";
endmodule

module DELAYA(A, LOAD_N, MOVE, DIRECTION, COARSE0, COARSE1, Z, EDETERR, CFLAG, RANKSELECT, RANKENABLE, RANK0UPDATE, RANK1UPDATE); //synthesis syn_black_box syn_lib_cell=1
    input A;
    input LOAD_N;
    input MOVE;
    input DIRECTION;
    input COARSE0;
    input COARSE1;
    input RANKSELECT;
    input RANKENABLE;
    input RANK0UPDATE;
    input RANK1UPDATE;
    output Z;
    output EDETERR;
    output CFLAG;
    parameter DEL_MODE = "USER_DEFINED";
    parameter DEL_VALUE = "0";
    parameter COARSE_DELAY_MODE = "STATIC";
    parameter COARSE_DELAY = "0NS";
    parameter EDGE_MONITOR = "DISABLED";
    parameter WAIT_FOR_EDGE = "DISABLED";
endmodule

module DELAYB(A, Z); //synthesis syn_black_box syn_lib_cell=1
    input A;
    output Z;
    parameter DEL_VALUE = "0";
    parameter COARSE_DELAY = "0NS";
    parameter DEL_MODE = "USER_DEFINED";
endmodule

module DELAYC(A, LOAD_N, MOVE, DIRECTION, COARSE0, COARSE1, Z, EDETERR, CFLAG, RANKSELECT, RANKENABLE, RANK0UPDATE, RANK1UPDATE, SCLK, ECLK); //synthesis syn_black_box syn_lib_cell=1
    input A;
    input LOAD_N;
    input MOVE; 
    input DIRECTION;
    input COARSE0;
    input COARSE1;
    output Z;
    output EDETERR;
    output CFLAG;
    input RANKSELECT;
    input RANKENABLE;
    input RANK0UPDATE;
    input RANK1UPDATE;
    input SCLK; 
    input ECLK; 
    parameter DEL_MODE = "USER_DEFINED";
    parameter DEL_VALUE = "0";
    parameter COARSE_DELAY_MODE = "STATIC";
    parameter COARSE_DELAY = "0NS";
    parameter EDGE_MONITOR = "DISABLED";
    parameter WAIT_FOR_EDGE = "DISABLED";
endmodule

module DIFFIO18(PADDO, DOLP, IOPAD, PADDI, INLP, PADDT, INADC, HSRXEN, HSTXEN); //synthesis black_box_pad_pin="IOPAD" syn_lib_cell=1
    input PADDO;
    input DOLP;
    inout IOPAD;
    output PADDI;
    output INLP;
    input PADDT;
    output INADC;
    input HSRXEN;
    input HSTXEN;
    parameter PULLMODE = "DOWN";
    parameter ENADC_IN = "DISABLED";
    parameter MIPI = "DISABLED";
endmodule

module DLLDEL(CLKIN, CLKOUT, CODE, COUT, DIR, LOAD_N, MOVE); //synthesis syn_black_box syn_lib_cell=1
    input CLKIN;
    output CLKOUT;
    input [8:0] CODE;
    output COUT;
    input DIR;
    input LOAD_N;
    input MOVE;
    parameter ADJUST = "0";
    parameter DEL_ADJUST = "PLUS";
    parameter ENABLE = "ENABLED";
endmodule

module DP16K_MODE(DIA0, DIA1, DIA2, DIA3, DIA4, DIA5, DIA6, DIA7, DIA8, DIA9, DIA10, DIA11, DIA12, DIA13, DIA14, DIA15, DIA16, DIA17, DIB0, DIB1, DIB2, DIB3, DIB4, DIB5, DIB6, DIB7, DIB8, DIB9, DIB10, DIB11, DIB12, DIB13, DIB14, DIB15, DIB16, DIB17, ADA0, ADA1, ADA2, ADA3, ADA4, ADA5, ADA6, ADA7, ADA8, ADA9, ADA10, ADA11, ADA12, ADA13, ADB0, ADB1, ADB2, ADB3, ADB4, ADB5, ADB6, ADB7, ADB8, ADB9, ADB10, ADB11, ADB12, ADB13, CLKA, CLKB, CEA, CEB, WEA, WEB, CSA0, CSA1, CSA2, CSB0, CSB1, CSB2, RSTA, RSTB, DOA0, DOA1, DOA2, DOA3, DOA4, DOA5, DOA6, DOA7, DOA8, DOA9, DOA10, DOA11, DOA12, DOA13, DOA14, DOA15, DOA16, DOA17, DOB0, DOB1, DOB2, DOB3, DOB4, DOB5, DOB6, DOB7, DOB8, DOB9, DOB10, DOB11, DOB12, DOB13, DOB14, DOB15, DOB16, DOB17); //synthesis syn_black_box syn_lib_cell=1
    input DIA0;
    input DIA1;
    input DIA2;
    input DIA3;
    input DIA4;
    input DIA5;
    input DIA6;
    input DIA7;
    input DIA8;
    input DIA9;
    input DIA10;
    input DIA11;
    input DIA12;
    input DIA13;
    input DIA14;
    input DIA15;
    input DIA16;
    input DIA17;
    input DIB0;
    input DIB1;
    input DIB2;
    input DIB3;
    input DIB4;
    input DIB5;
    input DIB6;
    input DIB7;
    input DIB8;
    input DIB9;
    input DIB10;
    input DIB11;
    input DIB12;
    input DIB13;
    input DIB14;
    input DIB15;
    input DIB16;
    input DIB17;
    input ADA0;
    input ADA1;
    input ADA2;
    input ADA3;
    input ADA4;
    input ADA5;
    input ADA6;
    input ADA7;
    input ADA8;
    input ADA9;
    input ADA10;
    input ADA11;
    input ADA12;
    input ADA13;
    input ADB0;
    input ADB1;
    input ADB2;
    input ADB3;
    input ADB4;
    input ADB5;
    input ADB6;
    input ADB7;
    input ADB8;
    input ADB9;
    input ADB10;
    input ADB11;
    input ADB12;
    input ADB13;
    input CLKA;
    input CLKB;
    input CEA;
    input CEB;
    input WEA;
    input WEB;
    input CSA0;
    input CSA1;
    input CSA2;
    input CSB0;
    input CSB1;
    input CSB2;
    input RSTA;
    input RSTB;
    output DOA0;
    output DOA1;
    output DOA2;
    output DOA3;
    output DOA4;
    output DOA5;
    output DOA6;
    output DOA7;
    output DOA8;
    output DOA9;
    output DOA10;
    output DOA11;
    output DOA12;
    output DOA13;
    output DOA14;
    output DOA15;
    output DOA16;
    output DOA17;
    output DOB0;
    output DOB1;
    output DOB2;
    output DOB3;
    output DOB4;
    output DOB5;
    output DOB6;
    output DOB7;
    output DOB8;
    output DOB9;
    output DOB10;
    output DOB11;
    output DOB12;
    output DOB13;
    output DOB14;
    output DOB15;
    output DOB16;
    output DOB17;
    parameter DATA_WIDTH_A = "X18";
    parameter DATA_WIDTH_B = "X18";
    parameter OUTREG_A = "BYPASSED";
    parameter OUTREG_B = "BYPASSED";
    parameter GSR = "ENABLED";
    parameter RESETMODE_A = "SYNC";
    parameter RESETMODE_B = "SYNC";
    parameter INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter CSDECODE_A = "000";
    parameter CSDECODE_B = "000";
    parameter ASYNC_RST_RELEASE_A = "SYNC";
    parameter ASYNC_RST_RELEASE_B = "SYNC";
    parameter INIT_DATA = "STATIC";
endmodule

module DP16K(DIA, DIB, ADA, ADB, CLKA, CLKB, CEA, CEB, WEA, WEB, CSA, CSB, RSTA, RSTB, DOA, DOB); //synthesis syn_black_box syn_lib_cell=1
    input [17:0] DIA;
    input [17:0] DIB;
    input [13:0] ADA;
    input [13:0] ADB;
    input CLKA;
    input CLKB;
    input CEA;
    input CEB;
    input WEA;
    input WEB;
    input [2:0] CSA;
    input [2:0] CSB;
    input RSTA;
    input RSTB;
    output [17:0] DOA;
    output [17:0] DOB;
    parameter DATA_WIDTH_A = "X18";
    parameter DATA_WIDTH_B = "X18";
    parameter OUTREG_A = "BYPASSED";
    parameter OUTREG_B = "BYPASSED";
    parameter GSR = "ENABLED";
    parameter RESETMODE_A = "SYNC";
    parameter RESETMODE_B = "SYNC";
    parameter INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter CSDECODE_A = "000";
    parameter CSDECODE_B = "000";
    parameter ASYNC_RST_RELEASE_A = "SYNC";
    parameter ASYNC_RST_RELEASE_B = "SYNC";
    parameter INIT_DATA = "STATIC";
endmodule

module DPHY(LMMICLK, LMMIRESET_N, LMMIREQUEST, LMMIWRRD_N, LMMIOFFSET, LMMIWDATA, LMMIRDATA, LMMIRDATAVALID, LMMIREADY, BITCKEXT, CKN, CKP, CLKREF, D0ACTIVE, D0BYTCNT, D0ERRCNT, D0PASS, D0VALID, D1ACTIVE, D1BYTCNT, D1ERRCNT, D1PASS, D1VALID, D2ACTIVE, D2BYTCNT, D2ERRCNT, D2PASS, D2VALID, D3ACTIVE, D3BYTCNT, D3ERRCNT, D3PASS, D3VALID, DCTSTOUT, DN0, DN1, DN2, DN3, DP0, DP1, DP2, DP3, LOCK, PDDPHY, PDPLL, SCCLKIN, UDIR, UED0THEN, UERCLP0, UERCLP1, UERCTRL, UERE, UERSTHS, UERSSHS, UERSE, UFRXMODE, UTXMDTX, URXACTHS, URXCKE, URXCKINE, URXDE, URXDHS, URXLPDTE, URXSKCHS, URXDRX, URXSHS, URE0D3DP, URE1D3DN, URE2CKDP, URE3CKDN, URXULPSE, URXVDE, URXVDHS, USSTT, UTDIS, UTXCKE, UDE0D0TN, UDE1D1TN, UDE2D2TN, UDE3D3TN, UDE4CKTN, UDE5D0RN, UDE6D1RN, UDE7D2RN, UTXDHS, UTXENER, UTXRRS, UTXRYP, UTXRYSK, UTXRD0EN, UTRD0SEN, UTXSKD0N, UTXTGE0, UTXTGE1, UTXTGE2, UTXTGE3, UTXULPSE, UTXUPSEX, UTXVDE, UTXWVDHS, UUSAN, U1DIR, U1ENTHEN, U1ERCLP0, U1ERCLP1, U1ERCTRL, U1ERE, U1ERSTHS, U1ERSSHS, U1ERSE, U1FRXMD, U1FTXST, U1RXATHS, U1RXCKE, U1RXDE, U1RXDHS, U1RXDTE, U1RXSKS, U1RXSK, U1RXSHS, U1RE0D, U1RE1CN, U1RE2D, U1RE3N, U1RXUPSE, U1RXVDE, U1RXVDHS, U1SSTT, U1TDIS, U1TREQ, U1TDE0D3, U1TDE1CK, U1TDE2D0, U1TDE3D1, U1TDE4D2, U1TDE5D3, U1TDE6, U1TDE7, U1TXDHS, U1TXLPD, U1TXRYE, U1TXRY, U1TXRYSK, U1TXREQ, U1TXREQH, U1TXSK, U1TXTGE0, U1TXTGE1, U1TXTGE2, U1TXTGE3, U1TXUPSE, U1TXUPSX, U1TXVDE, U1TXWVHS, U1USAN, U2DIR, U2END2, U2ERCLP0, U2ERCLP1, U2ERCTRL, U2ERE, U2ERSTHS, U2ERSSHS, U2ERSE, U2FRXMD, U2FTXST, U2RXACHS, U2RXCKE, U2RXDE, U2RXDHS, U2RPDTE, U2RXSK, U2RXSKC, U2RXSHS, U2RE0D2, U2RE1D2, U2RE2D3, U2RE3D3, U2RXUPSE, U2RXVDE, U2RXVDHS, U2SSTT, U2TDIS, U2TREQ, U2TDE0D0, U2TDE1D1, U2TDE2D2, U2TDE3D3, U2TDE4CK, U2TDE5D0, U2TDE6D1, U2TDE7D2, U2TXDHS, U2TPDTE, U2TXRYE, U2TXRYH, U2TXRYSK, U2TXREQ, U2TXREQH, U2TXSKC, U2TXTGE0, U2TXTGE1, U2TXTGE2, U2TXTGE3, U2TXUPSE, U2TXUPSX, U2TXVDE, U2TXWVHS, U2USAN, U3DIR, U3END3, U3ERCLP0, U3ERCLP1, U3ERCTRL, U3ERE, U3ERSTHS, U3ERSSHS, U3ERSE, U3FRXMD, U3FTXST, U3RXATHS, U3RXCKE, U3RXDE, U3RXDHS, U3RPDTE, U3RXSK, U3RXSKC, U3RXSHS, U3RE0CK, U3RE1CK, U3RE2, U3RE3, U3RXUPSE, U3RXVDE, U3RXVDHS, U3SSTT, U3TDISD2, U3TREQD2, U3TDE0D3, U3TDE1D0, U3TDE2D1, U3TDE3D2, U3TDE4D3, U3TDE5CK, U3TDE6, U3TDE7, U3TXDHS, U3TXLPDT, U3TXRY, U3TXRYHS, U3TXRYSK, U3TXREQ, U3TXREQH, U3TXSKC, U3TXTGE0, U3TXTGE1, U3TXTGE2, U3TXTGE3, U3TXULPS, U3TXUPSX, U3TXVD3, U3TXWVHS, U3USAN, UCENCK, UCRXCKAT, UCRXUCKN, UCSSTT, UCTXREQH, UCTXUPSC, UCTXUPSX, UCUSAN, LTSTEN, LTSTLANE, URWDCKHS, UTRNREQ, UTWDCKHS, UCRXWCHS, CLKLBACT); //synthesis black_box_pad_pin="CKN,CKP,DN0,DN1,DN2,DN3,DP0,DP1,DP2,DP3" syn_lib_cell=1
    input LMMICLK;
    input LMMIRESET_N;
    input LMMIREQUEST;
    input LMMIWRRD_N;
    input [4:0] LMMIOFFSET;
    input [3:0] LMMIWDATA;
    output [3:0] LMMIRDATA;
    output LMMIRDATAVALID;
    output LMMIREADY;
    input BITCKEXT;
    inout CKN;
    inout CKP;
    input CLKREF;
    output [1:0] D0ACTIVE;
    output [9:0] D0BYTCNT;
    output [9:0] D0ERRCNT;
    output [1:0] D0PASS;
    output [1:0] D0VALID;
    output [1:0] D1ACTIVE;
    output [9:0] D1BYTCNT;
    output [9:0] D1ERRCNT;
    output [1:0] D1PASS;
    output [1:0] D1VALID;
    output [1:0] D2ACTIVE;
    output [9:0] D2BYTCNT;
    output [9:0] D2ERRCNT;
    output [1:0] D2PASS;
    output [1:0] D2VALID;
    output [1:0] D3ACTIVE;
    output [9:0] D3BYTCNT;
    output [9:0] D3ERRCNT;
    output [1:0] D3PASS;
    output [1:0] D3VALID;
    output [9:0] DCTSTOUT;
    inout DN0;
    inout DN1;
    inout DN2;
    inout DN3;
    inout DP0;
    inout DP1;
    inout DP2;
    inout DP3;
    output LOCK;
    input PDDPHY;
    input PDPLL;
    input SCCLKIN;
    output UDIR;
    input UED0THEN;
    output UERCLP0;
    output UERCLP1;
    output UERCTRL;
    output UERE;
    output UERSTHS;
    output UERSSHS;
    output UERSE;
    input UFRXMODE;
    input UTXMDTX;
    output URXACTHS;
    output URXCKE;
    input URXCKINE;
    output [7:0] URXDE;
    output [15:0] URXDHS;
    output URXLPDTE;
    output URXSKCHS;
    output URXDRX;
    output [3:0] URXSHS;
    output URE0D3DP;
    output URE1D3DN;
    output URE2CKDP;
    output URE3CKDN;
    output URXULPSE;
    output URXVDE;
    output [3:0] URXVDHS;
    output USSTT;
    input UTDIS;
    input UTXCKE;
    input UDE0D0TN;
    input UDE1D1TN;
    input UDE2D2TN;
    input UDE3D3TN;
    input UDE4CKTN;
    input UDE5D0RN;
    input UDE6D1RN;
    input UDE7D2RN;
    input [31:0] UTXDHS;
    input UTXENER;
    output UTXRRS;
    output UTXRYP;
    output UTXRYSK;
    input UTXRD0EN;
    input UTRD0SEN;
    input UTXSKD0N;
    input UTXTGE0;
    input UTXTGE1;
    input UTXTGE2;
    input UTXTGE3;
    input UTXULPSE;
    input UTXUPSEX;
    input UTXVDE;
    input [3:0] UTXWVDHS;
    output UUSAN;
    output U1DIR;
    input U1ENTHEN;
    output U1ERCLP0;
    output U1ERCLP1;
    output U1ERCTRL;
    output U1ERE;
    output U1ERSTHS;
    output U1ERSSHS;
    output U1ERSE;
    input U1FRXMD;
    input U1FTXST;
    output U1RXATHS;
    output U1RXCKE;
    output [7:0] U1RXDE;
    output [15:0] U1RXDHS;
    output U1RXDTE;
    output U1RXSKS;
    output U1RXSK;
    output [3:0] U1RXSHS;
    output U1RE0D;
    output U1RE1CN;
    output U1RE2D;
    output U1RE3N;
    output U1RXUPSE;
    output U1RXVDE;
    output [3:0] U1RXVDHS;
    output U1SSTT;
    input U1TDIS;
    input U1TREQ;
    input U1TDE0D3;
    input U1TDE1CK;
    input U1TDE2D0;
    input U1TDE3D1;
    input U1TDE4D2;
    input U1TDE5D3;
    input U1TDE6;
    input U1TDE7;
    input [31:0] U1TXDHS;
    input U1TXLPD;
    output U1TXRYE;
    output U1TXRY;
    output U1TXRYSK;
    input U1TXREQ;
    input U1TXREQH;
    input U1TXSK;
    input U1TXTGE0;
    input U1TXTGE1;
    input U1TXTGE2;
    input U1TXTGE3;
    input U1TXUPSE;
    input U1TXUPSX;
    input U1TXVDE;
    input [3:0] U1TXWVHS;
    output U1USAN;
    output U2DIR;
    input U2END2;
    output U2ERCLP0;
    output U2ERCLP1;
    output U2ERCTRL;
    output U2ERE;
    output U2ERSTHS;
    output U2ERSSHS;
    output U2ERSE;
    input U2FRXMD;
    input U2FTXST;
    output U2RXACHS;
    output U2RXCKE;
    output [7:0] U2RXDE;
    output [15:0] U2RXDHS;
    output U2RPDTE;
    output U2RXSK;
    output U2RXSKC;
    output [3:0] U2RXSHS;
    output U2RE0D2;
    output U2RE1D2;
    output U2RE2D3;
    output U2RE3D3;
    output U2RXUPSE;
    output U2RXVDE;
    output [3:0] U2RXVDHS;
    output U2SSTT;
    input U2TDIS;
    input U2TREQ;
    input U2TDE0D0;
    input U2TDE1D1;
    input U2TDE2D2;
    input U2TDE3D3;
    input U2TDE4CK;
    input U2TDE5D0;
    input U2TDE6D1;
    input U2TDE7D2;
    input [31:0] U2TXDHS;
    input U2TPDTE;
    output U2TXRYE;
    output U2TXRYH;
    output U2TXRYSK;
    input U2TXREQ;
    input U2TXREQH;
    input U2TXSKC;
    input U2TXTGE0;
    input U2TXTGE1;
    input U2TXTGE2;
    input U2TXTGE3;
    input U2TXUPSE;
    input U2TXUPSX;
    input U2TXVDE;
    input [3:0] U2TXWVHS;
    output U2USAN;
    output U3DIR;
    input U3END3;
    output U3ERCLP0;
    output U3ERCLP1;
    output U3ERCTRL;
    output U3ERE;
    output U3ERSTHS;
    output U3ERSSHS;
    output U3ERSE;
    input U3FRXMD;
    input U3FTXST;
    output U3RXATHS;
    output U3RXCKE;
    output [7:0] U3RXDE;
    output [15:0] U3RXDHS;
    output U3RPDTE;
    output U3RXSK;
    output U3RXSKC;
    output [3:0] U3RXSHS;
    output U3RE0CK;
    output U3RE1CK;
    output U3RE2;
    output U3RE3;
    output U3RXUPSE;
    output U3RXVDE;
    output [3:0] U3RXVDHS;
    output U3SSTT;
    input U3TDISD2;
    input U3TREQD2;
    input U3TDE0D3;
    input U3TDE1D0;
    input U3TDE2D1;
    input U3TDE3D2;
    input U3TDE4D3;
    input U3TDE5CK;
    input U3TDE6;
    input U3TDE7;
    input [31:0] U3TXDHS;
    input U3TXLPDT;
    output U3TXRY;
    output U3TXRYHS;
    output U3TXRYSK;
    input U3TXREQ;
    input U3TXREQH;
    input U3TXSKC;
    input U3TXTGE0;
    input U3TXTGE1;
    input U3TXTGE2;
    input U3TXTGE3;
    input U3TXULPS;
    input U3TXUPSX;
    input U3TXVD3;
    input [3:0] U3TXWVHS;
    output U3USAN;
    input UCENCK;
    output UCRXCKAT;
    output UCRXUCKN;
    output UCSSTT;
    input UCTXREQH;
    input UCTXUPSC;
    input UCTXUPSX;
    output UCUSAN;
    input LTSTEN;
    input [1:0] LTSTLANE;
    output URWDCKHS;
    input UTRNREQ;
    output UTWDCKHS;
    output UCRXWCHS;
    output CLKLBACT;
    parameter GSR = "ENABLED";
    parameter AUTO_PD_EN = "POWERED_UP";
    parameter CFG_NUM_LANES = "ONE_LANE";
    parameter CM = "0b00000000";
    parameter CN = "0b00000";
    parameter CO = "0b000";
    parameter CONT_CLK_MODE = "DISABLED";
    parameter DESKEW_EN = "DISABLED";
    parameter DSI_CSI = "CSI2_APP";
    parameter EN_CIL = "CIL_ENABLED";
    parameter HSEL = "DISABLED";
    parameter LANE0_SEL = "LANE_0";
    parameter LOCK_BYP = "GATE_TXBYTECLKHS";
    parameter MASTER_SLAVE = "SLAVE";
    parameter PLLCLKBYPASS = "REGISTERED";
    parameter RSEL = "0b00";
    parameter RXCDRP = "0b00";
    parameter RXDATAWIDTHHS = "0b00";
    parameter RXLPRP = "0b000";
    parameter TEST_ENBL = "0b000000";
    parameter TEST_PATTERN = "0b00000000000000000000000000000000";
    parameter TST = "0b1001";
    parameter TXDATAWIDTHHS = "0b00";
    parameter U_PRG_HS_PREPARE = "0b00";
    parameter U_PRG_HS_TRAIL = "0b000000";
    parameter U_PRG_HS_ZERO = "0b000000";
    parameter U_PRG_RXHS_SETTLE = "0b000000";
    parameter UC_PRG_HS_PREPARE = "1P0_TXCLKESC";
    parameter UC_PRG_HS_TRAIL = "0b00000";
    parameter UC_PRG_HS_ZERO = "0b0000000";
    parameter UC_PRG_RXHS_SETTLE = "0b000000";
endmodule

module DPSC512K(DIA, DIB, ADA, ADB, CLK, CEA, CEB, WEA, WEB, CSA, CSB, RSTA, RSTB, BENA_N, BENB_N, CEOUTA, CEOUTB, DOA, DOB, ERRDECA, ERRDECB); //synthesis syn_black_box syn_lib_cell=1
    input [31:0] DIA;
    input [31:0] DIB;
    input [13:0] ADA;
    input [13:0] ADB;
    input CLK;
    input CEA;
    input CEB;
    input WEA;
    input WEB;
    input CSA;
    input CSB;
    input RSTA;
    input RSTB;
    input [3:0] BENA_N;
    input [3:0] BENB_N;
    input CEOUTA;
    input CEOUTB;
    output [31:0] DOA;
    output [31:0] DOB;
    output [1:0] ERRDECA;
    output [1:0] ERRDECB;
    parameter OUTREG_A = "NO_REG";
    parameter OUTREG_B = "NO_REG";
    parameter GSR = "ENABLED";
    parameter RESETMODE = "SYNC";
    parameter INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_40 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_41 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_42 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_43 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_44 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_45 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_46 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_47 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_48 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_49 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_4A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_4B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_4C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_4D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_4E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_4F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_50 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_51 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_52 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_53 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_54 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_55 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_56 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_57 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_58 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_59 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_5A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_5B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_5C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_5D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_5E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_5F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_60 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_61 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_62 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_63 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_64 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_65 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_66 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_67 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_68 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_69 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_6A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_6B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_6C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_6D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_6E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_6F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_70 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_71 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_72 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_73 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_74 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_75 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_76 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_77 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_78 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_79 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_7A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_7B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_7C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_7D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_7E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_7F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter ASYNC_RESET_RELEASE = "SYNC";
    parameter ECC_BYTE_SEL = "ECC_EN";
endmodule

module DQSBUF(BTDETECT, BURSTDETECT, DATAVALID, DQSI, DQSW, DQSWRD, PAUSE, RDCLKSEL, RDDIR, RDLOADN, RDPNTR, READ, READCOUT, READMOVE, RST, SCLK, SELCLK, DQSR90, DQSW270, WRCOUT, WRDIR, WRLOAD_N, WRLVCOUT, WRLVDIR, WRLVLOAD_N, WRLVMOVE, WRMOVE, WRPNTR, ECLKIN, RSTSMCNT, DLLCODE); //synthesis syn_black_box syn_lib_cell=1
    output BTDETECT;
    output BURSTDETECT;
    output DATAVALID;
    input DQSI;
    output DQSW;
    output DQSWRD;
    input PAUSE;
    input [3:0] RDCLKSEL;
    input RDDIR;
    input RDLOADN;
    output [2:0] RDPNTR;
    input [3:0] READ;
    output READCOUT;
    input READMOVE;
    input RST;
    input SCLK;
    input SELCLK;
    output DQSR90;
    output DQSW270;
    output WRCOUT;
    input WRDIR;
    input WRLOAD_N;
    output WRLVCOUT;
    input WRLVDIR;
    input WRLVLOAD_N;
    input WRLVMOVE;
    input WRMOVE;
    output [2:0] WRPNTR;
    input ECLKIN;
    input RSTSMCNT;
    input [8:0] DLLCODE;
    parameter GSR = "ENABLED";
    parameter ENABLE_FIFO = "DISABLED";
    parameter FORCE_READ = "DISABLED";
    parameter FREE_WHEEL = "DDR";
    parameter MODX = "NOT_USED";
    parameter MT_EN_READ = "DISABLED";
    parameter MT_EN_WRITE = "DISABLED";
    parameter MT_EN_WRITE_LEVELING = "DISABLED";
    parameter RD_PNTR = "0b000";
    parameter READ_ENABLE = "DISABLED";
    parameter RX_CENTERED = "ENABLED";
    parameter S_READ = "0";
    parameter S_WRITE = "0";
    parameter SIGN_READ = "POSITIVE";
    parameter SIGN_WRITE = "POSITIVE";
    parameter UPDATE_QU = "UP1_AND_UP0_SAME";
    parameter WRITE_ENABLE = "DISABLED";
    parameter SEL_READ_BIT_ENABLE_CYCLES = "NORMAL";
    parameter BYPASS_WR_LEVEL_SMTH_LATCH = "SMOOTHING_PATH";
    parameter BYPASS_WR_SMTH_LATCH = "SMOOTHING_PATH";
    parameter BYPASS_READ_SMTH_LATCH = "SMOOTHING_PATH";
endmodule

module EBR_CORE(DIA0, DIA1, DIA2, DIA3, DIA4, DIA5, DIA6, DIA7, DIA8, DIA9, DIA10, DIA11, DIA12, DIA13, DIA14, DIA15, DIA16, DIA17, DIB0, DIB1, DIB2, DIB3, DIB4, DIB5, DIB6, DIB7, DIB8, DIB9, DIB10, DIB11, DIB12, DIB13, DIB14, DIB15, DIB16, DIB17, ADA0, ADA1, ADA2, ADA3, ADA4, ADA5, ADA6, ADA7, ADA8, ADA9, ADA10, ADA11, ADA12, ADA13, ADB0, ADB1, ADB2, ADB3, ADB4, ADB5, ADB6, ADB7, ADB8, ADB9, ADB10, ADB11, ADB12, ADB13, CLKA, CLKB, WEA, WEB, CEA, CEB, RSTA, RSTB, CSA0, CSA1, CSA2, CSB0, CSB1, CSB2, FULLF, AFULL, EMPTYF, AEMPTY, DOA0, DOA1, DOA2, DOA3, DOA4, DOA5, DOA6, DOA7, DOA8, DOA9, DOA10, DOA11, DOA12, DOA13, DOA14, DOA15, DOA16, DOA17, DOB0, DOB1, DOB2, DOB3, DOB4, DOB5, DOB6, DOB7, DOB8, DOB9, DOB10, DOB11, DOB12, DOB13, DOB14, DOB15, DOB16, DOB17, ONEERR, TWOERR); //synthesis syn_black_box syn_lib_cell=1
    input DIA0;
    input DIA1;
    input DIA2;
    input DIA3;
    input DIA4;
    input DIA5;
    input DIA6;
    input DIA7;
    input DIA8;
    input DIA9;
    input DIA10;
    input DIA11;
    input DIA12;
    input DIA13;
    input DIA14;
    input DIA15;
    input DIA16;
    input DIA17;
    input DIB0;
    input DIB1;
    input DIB2;
    input DIB3;
    input DIB4;
    input DIB5;
    input DIB6;
    input DIB7;
    input DIB8;
    input DIB9;
    input DIB10;
    input DIB11;
    input DIB12;
    input DIB13;
    input DIB14;
    input DIB15;
    input DIB16;
    input DIB17;
    input ADA0;
    input ADA1;
    input ADA2;
    input ADA3;
    input ADA4;
    input ADA5;
    input ADA6;
    input ADA7;
    input ADA8;
    input ADA9;
    input ADA10;
    input ADA11;
    input ADA12;
    input ADA13;
    input ADB0;
    input ADB1;
    input ADB2;
    input ADB3;
    input ADB4;
    input ADB5;
    input ADB6;
    input ADB7;
    input ADB8;
    input ADB9;
    input ADB10;
    input ADB11;
    input ADB12;
    input ADB13;
    input CLKA;
    input CLKB;
    input WEA;
    input WEB;
    input CEA;
    input CEB;
    input RSTA;
    input RSTB;
    input CSA0;
    input CSA1;
    input CSA2;
    input CSB0;
    input CSB1;
    input CSB2;
    output FULLF;
    output AFULL;
    output EMPTYF;
    output AEMPTY;
    output DOA0;
    output DOA1;
    output DOA2;
    output DOA3;
    output DOA4;
    output DOA5;
    output DOA6;
    output DOA7;
    output DOA8;
    output DOA9;
    output DOA10;
    output DOA11;
    output DOA12;
    output DOA13;
    output DOA14;
    output DOA15;
    output DOA16;
    output DOA17;
    output DOB0;
    output DOB1;
    output DOB2;
    output DOB3;
    output DOB4;
    output DOB5;
    output DOB6;
    output DOB7;
    output DOB8;
    output DOB9;
    output DOB10;
    output DOB11;
    output DOB12;
    output DOB13;
    output DOB14;
    output DOB15;
    output DOB16;
    output DOB17;
    output ONEERR;
    output TWOERR;
    parameter INIT_DATA = "STATIC";
    parameter DATA_WIDTH_A = "X36";
    parameter DATA_WIDTH_B = "X36";
    parameter REGMODE_A = "BYPASSED";
    parameter REGMODE_B = "BYPASSED";
    parameter GSR = "ENABLED";
    parameter CSDECODE_A = "000";
    parameter CSDECODE_B = "000";
    parameter WID = "0b00000000000";
    parameter RESETMODE_A = "SYNC";
    parameter ASYNC_RESET_RELEASE_A = "SYNC";
    parameter RESETMODE_B = "SYNC";
    parameter ASYNC_RESET_RELEASE_B = "SYNC";
    parameter ECC = "DISABLED";
    parameter EBR_MODE = "DP";
    parameter FULL = "0b11111111100000";
    parameter ALMOST_FULL = "0b00000000000000";
    parameter EMPTY = "0b11111";
    parameter ALMOST_EMPTY = "0b00000000000000";
    parameter INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
endmodule

module EBR(DIA, DIB, ADA, ADB, CLKA, CLKB, WEA, WEB, CEA, CEB, RSTA, RSTB, CSA, CSB, FULLF, AFULL, EMPTYF, AEMPTY, DOA, DOB, ONEERR, TWOERR); //synthesis syn_black_box syn_lib_cell=1
    input [17:0] DIA;
    input [17:0] DIB;
    input [13:0] ADA;
    input [13:0] ADB;
    input CLKA;
    input CLKB;
    input WEA;
    input WEB;
    input CEA;
    input CEB;
    input RSTA;
    input RSTB;
    input [2:0] CSA;
    input [2:0] CSB;
    output FULLF;
    output AFULL;
    output EMPTYF;
    output AEMPTY;
    output [17:0] DOA;
    output [17:0] DOB;
    output ONEERR;
    output TWOERR;
    parameter INIT_DATA = "STATIC";
    parameter DATA_WIDTH_A = "X36";
    parameter DATA_WIDTH_B = "X36";
    parameter REGMODE_A = "BYPASSED";
    parameter REGMODE_B = "BYPASSED";
    parameter GSR = "ENABLED";
    parameter CSDECODE_A = "000";
    parameter CSDECODE_B = "000";
    parameter WID = "0b00000000000";
    parameter RESETMODE_A = "SYNC";
    parameter ASYNC_RESET_RELEASE_A = "SYNC";
    parameter RESETMODE_B = "SYNC";
    parameter ASYNC_RESET_RELEASE_B = "SYNC";
    parameter ECC = "DISABLED";
    parameter EBR_MODE = "DP";
    parameter FULL = "0b11111111100000";
    parameter ALMOST_FULL = "0b00000000000000";
    parameter ALMOST_EMPTY = "0b00000000000000";
    parameter INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
endmodule

module ECLKDIV(DIVOUT, DIVRST, ECLKIN, SLIP); //synthesis syn_black_box syn_lib_cell=1
    output DIVOUT;
    input DIVRST;
    input ECLKIN;
    input SLIP;
    parameter ECLK_DIV = "DISABLE";
    parameter GSR = "ENABLED";
endmodule

module ECLKSYNC(ECLKIN, ECLKOUT, STOP); //synthesis syn_black_box syn_lib_cell=1
    input ECLKIN;
    output ECLKOUT;
    input STOP;
    parameter STOP_EN = "DISABLE";
endmodule


module FBMUX(ENEXT, FBKCK, LGYRDYN, INTLOCK, WKUPSYNC, FBKCLK); //synthesis syn_black_box syn_lib_cell=1
    output ENEXT;
    output FBKCK;
    input LGYRDYN;
    input INTLOCK;
    input WKUPSYNC;
    input [15:0] FBKCLK;
    parameter INTFB = "IGNORED";
    parameter SEL_FBK = "DIVA";
    parameter CLKMUX_FB = "CMUX_CLKOP";
    parameter INTFBKDEL_SEL = "DISABLED";
endmodule


module FIFO16K_MODE(DI0, DI1, DI2, DI3, DI4, DI5, DI6, DI7, DI8, DI9, DI10,DI11, DI12, DI13, DI14, DI15, DI16, DI17, DI18, DI19, DI20,DI21, DI22, DI23, DI24, DI25, DI26, DI27, DI28, DI29, DI30,DI31, DI32, DI33, DI34, DI35,CLKW, CLKR,WE, RE,RSTW, RPRST,FULLI, EMPTYI,CSW0, CSW1,CSR0, CSR1,DO0, DO1, DO2, DO3, DO4, DO5, DO6, DO7, DO8, DO9, DO10,DO11, DO12, DO13, DO14, DO15, DO16, DO17, DO18, DO19, DO20,DO21, DO22, DO23, DO24, DO25, DO26, DO27, DO28, DO29, DO30,DO31, DO32, DO33, DO34, DO35,ONEBITERR, TWOBITERR,ALMOSTFULL, FULL, ALMOSTEMPTY, EMPTY); //synthesis syn_black_box syn_lib_cell=1
    input DI0;
    input DI1;
    input DI2;
    input DI3;
    input DI4;
    input DI5;
    input DI6;
    input DI7;
    input DI8;
    input DI9;
    input DI10;
    input DI11;
    input DI12;
    input DI13;
    input DI14;
    input DI15;
    input DI16;
    input DI17;
    input DI18;
    input DI19;
    input DI20;
    input DI21;
    input DI22;
    input DI23;
    input DI24;
    input DI25;
    input DI26;
    input DI27;
    input DI28;
    input DI29;
    input DI30;
    input DI31;
    input DI32;
    input DI33;
    input DI34;
    input DI35;
    input CLKW;
    input CLKR;
    input WE;
    input RE;
    input RSTW;
    input RPRST;
    input FULLI;
    input EMPTYI;
    input CSW0;
    input CSW1;
    input CSR0;
    input CSR1;
    output DO0;
    output DO1;
    output DO2;
    output DO3;
    output DO4;
    output DO5;
    output DO6;
    output DO7;
    output DO8;
    output DO9;
    output DO10;
    output DO11;
    output DO12;
    output DO13;
    output DO14;
    output DO15;
    output DO16;
    output DO17;
    output DO18;
    output DO19;
    output DO20;
    output DO21;
    output DO22;
    output DO23;
    output DO24;
    output DO25;
    output DO26;
    output DO27;
    output DO28;
    output DO29;
    output DO30;
    output DO31;
    output DO32;
    output DO33;
    output DO34;
    output DO35;
    output ONEBITERR;
    output TWOBITERR;
    output ALMOSTFULL;
    output FULL;
    output ALMOSTEMPTY;
    output EMPTY;
    parameter DATA_WIDTH_W = "X36";
    parameter DATA_WIDTH_R = "X36";
    parameter OUTREG = "BYPASSED";
    parameter GSR = "ENABLED";
    parameter RESETMODE = "SYNC";
    parameter ASYNC_RST_RELEASE = "SYNC";
    parameter ECC = "DISABLED";
    parameter CSDECODE_W = "00";
    parameter CSDECODE_R = "00";
    parameter FULLBITS = "0b10000000000000";
    parameter ALMOST_FULL = "0b00000000000000";
    parameter ALMOST_EMPTY = "0b00000000000000";
endmodule

module FIFO16K(DI, CLKW, CLKR, WE, RE, RSTW, RPRST, FULLI, EMPTYI, CSW, CSR, DO, ONEBITERR, TWOBITERR, ALMOSTFULL, FULL, ALMOSTEMPTY, EMPTY); //synthesis syn_black_box syn_lib_cell=1
    input [35:0] DI;
    input CLKW;
    input CLKR;
    input WE;
    input RE;
    input RSTW;
    input RPRST;
    input FULLI;
    input EMPTYI;
    input [1:0] CSW;
    input [1:0] CSR;
    output [35:0] DO;
    output ONEBITERR;
    output TWOBITERR;
    output ALMOSTFULL;
    output FULL;
    output ALMOSTEMPTY;
    output EMPTY;
    parameter DATA_WIDTH_W = "X36";
    parameter DATA_WIDTH_R = "X36";
    parameter OUTREG = "BYPASSED";
    parameter GSR = "ENABLED";
    parameter RESETMODE = "SYNC";
    parameter ASYNC_RST_RELEASE = "SYNC";
    parameter ECC = "DISABLED";
    parameter CSDECODE_W = "00";
    parameter CSDECODE_R = "00";
    parameter FULLBITS = "0b10000000000000";
    parameter ALMOST_FULL = "0b00000000000000";
    parameter ALMOST_EMPTY = "0b00000000000000";
endmodule

// R2.1 :
// module CRE taken out from je5d00/lifcl
// R2.2 : added back, will be stripped by relman build,
// & added to controlpack_cre during relman build.
//


module I2CFIFO(LMMICLK, LMMIRESET_N, LMMIREQUEST, LMMIWRRD_N, LMMIOFFSET, LMMIWDATA, LMMIRDATA, LMMIRDATAVALID, LMMIREADY, ALTSCLIN, ALTSCLOEN, ALTSCLOUT, ALTSDAIN, ALTSDAOEN, ALTSDAOUT, BUSBUSY, FIFORESET, I2CLSRRSTN, INSLEEP, IRQ, MRDCMPL, RXFIFOAF, RXFIFOE, RXFIFOF, SCLIN, SCLOE, SCLOEN, SCLOUT, SDAIN, SDAOE, SDAOEN, SDAOUT, SLVADDRMATCH, SLVADDRMATCHSCL, SRDWR, TXFIFOAE, TXFIFOE, TXFIFOF); //synthesis syn_black_box syn_lib_cell=1
    input LMMICLK;
    input LMMIRESET_N;
    input LMMIREQUEST;
    input LMMIWRRD_N;
    input [5:0] LMMIOFFSET;
    input [7:0] LMMIWDATA;
    output [7:0] LMMIRDATA;
    output LMMIRDATAVALID;
    output LMMIREADY;
    input ALTSCLIN;
    output ALTSCLOEN;
    output ALTSCLOUT;
    input ALTSDAIN;
    output ALTSDAOEN;
    output ALTSDAOUT;
    output BUSBUSY;
    input FIFORESET;
    input I2CLSRRSTN;
    output INSLEEP;
    output IRQ;
    output MRDCMPL;
    output RXFIFOAF;
    output RXFIFOE;
    output RXFIFOF;
    input SCLIN;
    output SCLOE;
    output SCLOEN;
    output SCLOUT;
    input SDAIN;
    output SDAOE;
    output SDAOEN;
    output SDAOUT;
    output SLVADDRMATCH;
    output SLVADDRMATCHSCL;
    output SRDWR;
    output TXFIFOAE;
    output TXFIFOE;
    output TXFIFOF;
    parameter BRNBASEDELAY = "0b0000";
    parameter CR1CKDIS = "EN";
    parameter CR1FIFOMODE = "REG";
    parameter CR1GCEN = "DIS";
    parameter CR1I2CEN = "DIS";
    parameter CR1SDADELSEL = "NDLY0";
    parameter CR1SLPCLKEN = "DIS";
    parameter CR2CORERSTN = "DIS";
    parameter CR2HARDTIE = "TIE";
    parameter CR2INTCLREN = "DIS";
    parameter CR2MRDCMPLWKUP = "DIS";
    parameter CR2RXFIFOAFWKUP = "DIS";
    parameter CR2SLVADDRWKUP = "DIS";
    parameter GSR = "ENABLED";
    parameter I2CADDRSEL = "7BIT";
    parameter I2CRXFIFOAFVAL = "0b00000";
    parameter I2CSLVADDRA = "0b0000000000";
    parameter I2CTXFIFOAEVAL = "0b0000";
    parameter INTARBLIE = "DIS";
    parameter INTBUSFREEIE = "DIS";
    parameter INTHGCIE = "DIS";
    parameter INTMRDCMPLIE = "DIS";
    parameter INTRNACKIEORRSVD = "DIS";
    parameter INTRSVDORTROEIE = "DIS";
    parameter INTRSVDORTRRDYIE = "DIS";
    parameter INTRXOVERFIEORRSVD = "DIS";
    parameter INTRXUNDERFIE = "DIS";
    parameter INTTXOVERFIE = "DIS";
    parameter INTTXSERRIEORRSVD = "DIS";
    parameter LMMI_EXTRA_ONE = "DIS";
    parameter LMMI_EXTRA_TWO = "DIS";
    parameter NCRALTIOEN = "FABRIC";
    parameter NCRFILTERDIS = "EN";
    parameter NCRSDAINDLYEN = "DIS";
    parameter NCRSDAOUTDLYEN = "DIS";
    parameter NONUSRTESTSOFTTRIMEN = "DIS";
    parameter NONUSRTSTSOFTTRIMVALUE = "0b000";
    parameter REGI2CBR = "0b0000000000";
    parameter TSPTIMERVALUE = "0b10010010111";
endmodule

module IDDR71(D, SCLK, RST, ECLK, ALIGNWD, Q0, Q1, Q2, Q3, Q4, Q5, Q6); //synthesis syn_black_box syn_lib_cell=1
    input D;
    input SCLK;
    input RST;
    input ECLK;
    input ALIGNWD;
    output Q0;
    output Q1;
    output Q2;
    output Q3;
    output Q4;
    output Q5;
    output Q6;
    parameter GSR = "ENABLED";
endmodule

module IDDRX1(D, SCLK, RST, Q0, Q1); //synthesis syn_black_box syn_lib_cell=1
    input D;
    input SCLK;
    input RST;
    output Q0;
    output Q1;
    parameter GSR = "ENABLED";
endmodule

module IDDRX2DQ(D, DQSR90, ECLK, SCLK, RST, RDPNTR0, RDPNTR1, RDPNTR2, WRPNTR0, WRPNTR1, WRPNTR2, Q0, Q1, Q2, Q3); //synthesis syn_black_box syn_lib_cell=1
    input D;
    input DQSR90;
    input ECLK;
    input SCLK;
    input RST;
    input RDPNTR0;
    input RDPNTR1;
    input RDPNTR2;
    input WRPNTR0;
    input WRPNTR1;
    input WRPNTR2;
    output Q0;
    output Q1;
    output Q2;
    output Q3;
    parameter GSR = "ENABLED";
endmodule

module IDDRX2(D, SCLK, RST, ECLK, ALIGNWD, Q0, Q1, Q2, Q3); //synthesis syn_black_box syn_lib_cell=1
    input D;
    input SCLK;
    input RST;
    input ECLK;
    input ALIGNWD;
    output Q0;
    output Q1;
    output Q2;
    output Q3;
    parameter GSR = "ENABLED";
endmodule

module IDDRX4DQ(D, DQSR90, ECLK, SCLK, RST, RDPNTR0, RDPNTR1, RDPNTR2, WRPNTR0, WRPNTR1, WRPNTR2, Q0, Q1, Q2, Q3, Q4, Q5, Q6, Q7); //synthesis syn_black_box syn_lib_cell=1
    input D;
    input DQSR90;
    input ECLK;
    input SCLK;
    input RST;
    input RDPNTR0;
    input RDPNTR1;
    input RDPNTR2;
    input WRPNTR0;
    input WRPNTR1;
    input WRPNTR2;
    output Q0;
    output Q1;
    output Q2;
    output Q3;
    output Q4;
    output Q5;
    output Q6;
    output Q7;
    parameter GSR = "ENABLED";
endmodule

module IDDRX4(D, SCLK, RST, ECLK, ALIGNWD, Q0, Q1, Q2, Q3, Q4, Q5, Q6, Q7); //synthesis syn_black_box syn_lib_cell=1
    input D;
    input SCLK;
    input RST;
    input ECLK;
    input ALIGNWD;
    output Q0;
    output Q1;
    output Q2;
    output Q3;
    output Q4;
    output Q5;
    output Q6;
    output Q7;
    parameter GSR = "ENABLED";
endmodule

module IDDRX5(D, SCLK, RST, ECLK, ALIGNWD, Q0, Q1, Q2, Q3, Q4, Q5, Q6, Q7, Q8, Q9); //synthesis syn_black_box syn_lib_cell=1
    input D;
    input SCLK;
    input RST;
    input ECLK;
    input ALIGNWD;
    output Q0;
    output Q1;
    output Q2;
    output Q3;
    output Q4;
    output Q5;
    output Q6;
    output Q7;
    output Q8;
    output Q9;
    parameter GSR = "ENABLED";
endmodule

module IFD1P3BX(D, SP, CK, PD, Q); //synthesis syn_black_box syn_lib_cell=1
    input D;
    input SP;
    input CK;
    input PD;
    output Q;
    parameter GSR = "ENABLED";
endmodule

module IFD1P3DX(D, SP, CK, CD, Q); //synthesis syn_black_box syn_lib_cell=1
    input D;
    input SP;
    input CK;
    input CD;
    output Q;
    parameter GSR = "ENABLED";
endmodule

module IFD1P3IX(D, SP, CK, CD, Q); //synthesis syn_black_box syn_lib_cell=1
    input D;
    input SP;
    input CK;
    input CD;
    output Q;
    parameter GSR = "ENABLED";
endmodule

module IFD1P3JX(D, SP, CK, PD, Q); //synthesis syn_black_box syn_lib_cell=1
    input D;
    input SP;
    input CK;
    input PD;
    output Q;
    parameter GSR = "ENABLED";
endmodule

module JTAG(JCE1, JCE2, JRSTN, JRTI1, JRTI2, JSHIFT, JTDI, JUPDATE, JTDO1, JTDO2, SMCLK, TCK, JTCK, TDI, TDO_OEN, TDO, TMS); //synthesis syn_black_box syn_lib_cell=1
    output JCE1;
    output JCE2;
    output JRSTN;
    output JRTI1;
    output JRTI2;
    output JSHIFT;
    output JTDI;
    output JUPDATE;
    input JTDO1;
    input JTDO2;
    input SMCLK;
    input TCK;
    output JTCK;
    input TDI;
    output TDO_OEN;
    output TDO;
    input TMS;
    parameter MCER1EXIST = "NEXIST";
    parameter MCER2EXIST = "NEXIST";
endmodule

module LRAM(ADA, ADB, BENA_N, BENB_N, CEA, CEB, CLK, CSA, CSB, DIA, DIB, DOA, DOB, DPS, ERRDECA, ERRDECB, OCEA, OCEB, OEA, OEB, RSTA, RSTB, WEA, WEB, ERRDET, LRAMREADY); //synthesis syn_black_box syn_lib_cell=1
    input [13:0] ADA;
    input [13:0] ADB;
    input [3:0] BENA_N;
    input [3:0] BENB_N;
    input CEA;
    input CEB;
    input CLK;
    input CSA;
    input CSB;
    input [31:0] DIA;
    input [31:0] DIB;
    output [31:0] DOA;
    output [31:0] DOB;
    input DPS;
    output [1:0] ERRDECA;
    output [1:0] ERRDECB;
    input OCEA;
    input OCEB;
    output OEA;
    output OEB;
    input RSTA;
    input RSTB;
    input WEA;
    input WEB;
    output ERRDET;
    output LRAMREADY;
    parameter INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_40 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_41 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_42 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_43 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_44 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_45 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_46 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_47 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_48 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_49 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_4A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_4B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_4C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_4D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_4E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_4F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_50 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_51 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_52 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_53 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_54 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_55 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_56 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_57 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_58 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_59 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_5A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_5B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_5C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_5D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_5E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_5F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_60 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_61 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_62 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_63 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_64 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_65 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_66 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_67 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_68 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_69 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_6A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_6B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_6C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_6D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_6E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_6F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_70 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_71 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_72 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_73 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_74 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_75 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_76 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_77 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_78 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_79 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_7A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_7B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_7C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_7D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_7E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_7F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter ASYNC_RST_RELEASE = "SYNC";
    parameter CFG_INIT_ID = "0b00000000000";
    parameter DATA_PRESERVE = "DISABLE";
    parameter EBR_SP_EN = "DISABLE";
    parameter ECC_BYTE_SEL = "ECC_EN";
    parameter GSR = "ENABLED";
    parameter OUT_REGMODE_A = "NO_REG";
    parameter OUT_REGMODE_B = "NO_REG";
    parameter RESETMODE = "SYNC";
    parameter RST_AB_EN = "RESET_AB_DISABLE";
    parameter SP_EN = "DISABLE";
    parameter UNALIGNED_READ = "DISABLE";
endmodule

module M18X36(SFTCTRL, PH36, PL36, SGNED18H, SGNED18L, P72, ROUNDEN); //synthesis syn_black_box syn_lib_cell=1
    input [3:0] SFTCTRL;
    input [37:0] PH36;
    input [37:0] PL36;
    input SGNED18H;
    input SGNED18L;
    output [72:0] P72;
    input ROUNDEN;
    parameter SFTEN = "DISABLED";
    parameter MULT18X36 = "ENABLED";
    parameter MULT36 = "DISABLED";
    parameter MULT36X36H = "USED_AS_LOWER_BIT_GENERATION";
    parameter ROUNDHALFUP = "DISABLED";
    parameter ROUNDRTZI = "ROUND_TO_ZERO";
    parameter ROUNDBIT = "ROUND_TO_BIT0";
endmodule

module MULT18(SFTCTRL, ARHSIGN, BRHSIGN, ARH, BRH, ARL, BRL, PL18, PH18, SIGNED18, P36, ROUNDEN); //synthesis syn_black_box syn_lib_cell=1
    input [3:0] SFTCTRL;
    input ARHSIGN;
    input BRHSIGN;
    input [8:0] ARH;
    input [8:0] BRH;
    input [8:0] ARL;
    input [8:0] BRL;
    input [19:0] PL18;
    input [19:0] PH18;
    output SIGNED18;
    output [37:0] P36;
    input ROUNDEN;
    parameter SFTEN = "DISABLED";
    parameter MULT18X18 = "ENABLED";
    parameter ROUNDHALFUP = "DISABLED";
    parameter ROUNDRTZI = "ROUND_TO_ZERO";
    parameter ROUNDBIT = "ROUND_TO_BIT0";
endmodule

module MULT18X18(A, B, CLK, CEA, RSTA, CEB, RSTB, SIGNEDA, SIGNEDB, RSTOUT, CEOUT, Z); //synthesis syn_black_box syn_lib_cell=1
    input [17:0] A;
    input [17:0] B;
    input CLK;
    input CEA;
    input RSTA;
    input CEB;
    input RSTB;
    input SIGNEDA;
    input SIGNEDB;
    input RSTOUT;
    input CEOUT;
    output [35:0] Z;
    parameter REGINPUTA = "REGISTER";
    parameter REGINPUTB = "REGISTER";
    parameter REGOUTPUT = "REGISTER";
    parameter GSR = "ENABLED";
    parameter RESETMODE = "SYNC";
endmodule

module MULT18X36(A, B, CLK, CEA, RSTA, CEB, RSTB, SIGNEDA, SIGNEDB, RSTOUT, CEOUT, Z); //synthesis syn_black_box syn_lib_cell=1
    input [17:0] A;
    input [35:0] B;
    input CLK;
    input CEA;
    input RSTA;
    input CEB;
    input RSTB;
    input SIGNEDA;
    input SIGNEDB;
    input RSTOUT;
    input CEOUT;
    output [53:0] Z;
    parameter REGINPUTA = "REGISTER";
    parameter REGINPUTB = "REGISTER";
    parameter REGOUTPUT = "REGISTER";
    parameter GSR = "ENABLED";
    parameter RESETMODE = "SYNC";
endmodule

module MULT36(PH72, PL72, PML72, PMH72); //synthesis syn_black_box syn_lib_cell=1
    input [72:0] PH72;
    input [72:0] PL72;
    output [71:0] PML72;
    output [71:0] PMH72;
    parameter MULT36X36 = "ENABLED";
endmodule

module MULT36X36(A, B, CLK, CEA, RSTA, CEB, RSTB, SIGNEDA, SIGNEDB, RSTOUT, CEOUT, Z); //synthesis syn_black_box syn_lib_cell=1
    input [35:0] A;
    input [35:0] B;
    input CLK;
    input CEA;
    input RSTA;
    input CEB;
    input RSTB;
    input SIGNEDA;
    input SIGNEDB;
    input RSTOUT;
    input CEOUT;
    output [71:0] Z;
    parameter REGINPUTA = "REGISTER";
    parameter REGINPUTB = "REGISTER";
    parameter REGOUTPUT = "REGISTER";
    parameter GSR = "ENABLED";
    parameter RESETMODE = "SYNC";
endmodule

module MULT9(A, ASIGNED, BR, AS1, AS2, ASSIGNED1, ASSIGNED2, BRSIGNED, CLK, CEA, RSTA, AO, BO, AOSIGNED, BOSIGNED, AR, ARSIGNED, P18, CEP, RSTP); //synthesis syn_black_box syn_lib_cell=1
    input [8:0] A;
    input ASIGNED;
    input [8:0] BR;
    input [8:0] AS1;
    input [8:0] AS2;
    input ASSIGNED1;
    input ASSIGNED2;
    input BRSIGNED;
    input CLK;
    input CEA;
    input RSTA;
    output [8:0] AO;
    output [8:0] BO;
    output AOSIGNED;
    output BOSIGNED;
    output [8:0] AR;
    output ARSIGNED;
    output [19:0] P18;
    input CEP;
    input RSTP;
    parameter SIGNEDSTATIC_EN = "DISABLED";
    parameter ASIGNED_OPERAND_EN = "DISABLED";
    parameter BYPASS_MULT9 = "USED";
    parameter REGBYPSB = "REGISTER";
    parameter REGBYPSA1 = "REGISTER";
    parameter REGBYPSA2 = "REGISTER";
    parameter SHIFTA = "DISABLED";
    parameter SR_18BITSHIFT_EN = "DISABLED";
    parameter GSR = "ENABLED";
    parameter RESET = "SYNC";
endmodule

module MULT9X9(A, B, CLK, CEA, RSTA, CEB, RSTB, SIGNEDA, SIGNEDB, RSTOUT, CEOUT, Z); //synthesis syn_black_box syn_lib_cell=1
    input [8:0] A;
    input [8:0] B;
    input CLK;
    input CEA;
    input RSTA;
    input CEB;
    input RSTB;
    input SIGNEDA;
    input SIGNEDB;
    input RSTOUT;
    input CEOUT;
    output [17:0] Z;
    parameter REGINPUTA = "REGISTER";
    parameter REGINPUTB = "REGISTER";
    parameter REGOUTPUT = "REGISTER";
    parameter GSR = "ENABLED";
    parameter RESETMODE = "SYNC";
endmodule

module MULTADDSUB18X18(A, B, C, CLK, CEA, RSTA, CEB, RSTB, CEC, RSTC, SIGNED, RSTPIPE, CEPIPE, RSTCTRL, CECTRL, RSTCIN, CECIN, LOADC, ADDSUB, Z, RSTOUT, CEOUT, CIN); //synthesis syn_black_box syn_lib_cell=1
    input [17:0] A;
    input [17:0] B;
    input [53:0] C;
    input CLK;
    input CEA;
    input RSTA;
    input CEB;
    input RSTB;
    input CEC;
    input RSTC;
    input SIGNED;
    input RSTPIPE;
    input CEPIPE;
    input RSTCTRL;
    input CECTRL;
    input RSTCIN;
    input CECIN;
    input LOADC;
    input ADDSUB;
    output [53:0] Z;
    input RSTOUT;
    input CEOUT;
    input CIN;
    parameter REGINPUTA = "REGISTER";
    parameter REGINPUTB = "REGISTER";
    parameter REGINPUTC = "REGISTER";
    parameter REGADDSUB = "REGISTER";
    parameter REGLOADC = "REGISTER";
    parameter REGLOADC2 = "REGISTER";
    parameter REGCIN = "REGISTER";
    parameter REGPIPELINE = "REGISTER";
    parameter REGOUTPUT = "REGISTER";
    parameter GSR = "ENABLED";
    parameter RESETMODE = "SYNC";
endmodule

module MULTADDSUB18X18WIDE(A0, B0, A1, B1, C, CLK, CEA0, CEA1, RSTA0, RSTA1, CEB0, CEB1, RSTB0, RSTB1, CEC, RSTC, RSTCTRL, CECTRL, SIGNED, RSTPIPE, CEPIPE, Z, RSTOUT, CEOUT, LOADC, ADDSUB); //synthesis syn_black_box syn_lib_cell=1
    input [17:0] A0;
    input [17:0] B0;
    input [17:0] A1;
    input [17:0] B1;
    input [53:0] C;
    input CLK;
    input CEA0;
    input CEA1;
    input RSTA0;
    input RSTA1;
    input CEB0;
    input CEB1;
    input RSTB0;
    input RSTB1;
    input CEC;
    input RSTC;
    input RSTCTRL;
    input CECTRL;
    input SIGNED;
    input RSTPIPE;
    input CEPIPE;
    output [53:0] Z;
    input RSTOUT;
    input CEOUT;
    input LOADC;
    input [1:0] ADDSUB;
    parameter REGINPUTAB0 = "REGISTER";
    parameter REGINPUTAB1 = "REGISTER";
    parameter REGINPUTC = "REGISTER";
    parameter REGADDSUB = "REGISTER";
    parameter REGLOADC = "REGISTER";
    parameter REGLOADC2 = "REGISTER";
    parameter REGPIPELINE = "REGISTER";
    parameter REGOUTPUT = "REGISTER";
    parameter GSR = "ENABLED";
    parameter RESETMODE = "SYNC";
endmodule

module MULTADDSUB18X36(A, B, C, CLK, CEA, RSTA, CEB, RSTB, CEC, RSTC, RSTCTRL, CECTRL, RSTCIN, CECIN, SIGNED, RSTPIPE, CEPIPE, RSTOUT, CEOUT, Z, LOADC, ADDSUB, CIN); //synthesis syn_black_box syn_lib_cell=1
    input [17:0] A;
    input [35:0] B;
    input [53:0] C;
    input CLK;
    input CEA;
    input RSTA;
    input CEB;
    input RSTB;
    input CEC;
    input RSTC;
    input RSTCTRL;
    input CECTRL;
    input RSTCIN;
    input CECIN;
    input SIGNED;
    input RSTPIPE;
    input CEPIPE;
    input RSTOUT;
    input CEOUT;
    output [53:0] Z;
    input LOADC;
    input ADDSUB;
    input CIN;
    parameter REGINPUTA = "REGISTER";
    parameter REGINPUTB = "REGISTER";
    parameter REGINPUTC = "REGISTER";
    parameter REGADDSUB = "REGISTER";
    parameter REGLOADC = "REGISTER";
    parameter REGLOADC2 = "REGISTER";
    parameter REGCIN = "REGISTER";
    parameter REGPIPELINE = "REGISTER";
    parameter REGOUTPUT = "REGISTER";
    parameter GSR = "ENABLED";
    parameter RESETMODE = "SYNC";
endmodule

module MULTADDSUB36X36(A, B, C, CLK, CEA, RSTA, CEB, RSTB, CEC, RSTC, RSTCTRL, CECTRL, RSTCIN, CECIN, SIGNED, RSTPIPE, CEPIPE, RSTOUT, CEOUT, Z, LOADC, ADDSUB, CIN); //synthesis syn_black_box syn_lib_cell=1
    input [35:0] A;
    input [35:0] B;
    input [107:0] C;
    input CLK;
    input CEA;
    input RSTA;
    input CEB;
    input RSTB;
    input CEC;
    input RSTC;
    input RSTCTRL;
    input CECTRL;
    input RSTCIN;
    input CECIN;
    input SIGNED;
    input RSTPIPE;
    input CEPIPE;
    input RSTOUT;
    input CEOUT;
    output [107:0] Z;
    input LOADC;
    input ADDSUB;
    input CIN;
    parameter REGINPUTA = "REGISTER";
    parameter REGINPUTB = "REGISTER";
    parameter REGINPUTC = "REGISTER";
    parameter REGADDSUB = "REGISTER";
    parameter REGLOADC = "REGISTER";
    parameter REGLOADC2 = "REGISTER";
    parameter REGCIN = "REGISTER";
    parameter REGPIPELINE = "REGISTER";
    parameter REGOUTPUT = "REGISTER";
    parameter GSR = "ENABLED";
    parameter RESETMODE = "SYNC";
endmodule

module MULTADDSUB9X9WIDE(A0, B0, A1, B1, A2, B2, A3, B3, C, CLK, CEA0A1, CEA2A3, RSTA0A1, RSTA2A3, CEB0B1, CEB2B3, RSTB0B1, RSTB2B3, CEC, RSTC, RSTCTRL, CECTRL, SIGNED, RSTPIPE, CEPIPE, RSTOUT, CEOUT, LOADC, ADDSUB, Z); //synthesis syn_black_box syn_lib_cell=1
    input [8:0] A0;
    input [8:0] B0;
    input [8:0] A1;
    input [8:0] B1;
    input [8:0] A2;
    input [8:0] B2;
    input [8:0] A3;
    input [8:0] B3;
    input [53:0] C;
    input CLK;
    input CEA0A1;
    input CEA2A3;
    input RSTA0A1;
    input RSTA2A3;
    input CEB0B1;
    input CEB2B3;
    input RSTB0B1;
    input RSTB2B3;
    input CEC;
    input RSTC;
    input RSTCTRL;
    input CECTRL;
    input SIGNED;
    input RSTPIPE;
    input CEPIPE;
    input RSTOUT;
    input CEOUT;
    input LOADC;
    input [3:0] ADDSUB;
    output [53:0] Z;
    parameter REGINPUTAB0 = "REGISTER";
    parameter REGINPUTAB1 = "REGISTER";
    parameter REGINPUTAB2 = "REGISTER";
    parameter REGINPUTAB3 = "REGISTER";
    parameter REGINPUTC = "REGISTER";
    parameter REGADDSUB = "REGISTER";
    parameter REGLOADC = "REGISTER";
    parameter REGLOADC2 = "REGISTER";
    parameter REGPIPELINE = "REGISTER";
    parameter REGOUTPUT = "REGISTER";
    parameter GSR = "ENABLED";
    parameter RESETMODE = "SYNC";
endmodule

module MULTIBOOT(AUTOREBOOT, MSPIMADDR); //synthesis syn_noprune=1 syn_lib_cell=1
    input AUTOREBOOT;
    input [31:0] MSPIMADDR;
    parameter MSPIADDR = "0b00000000000000000000000000000000";
    parameter SOURCESEL = "DIS";
endmodule

module MULTPREADD18X18(A, B, C, CLK, CEA, RSTA, CEB, RSTB, CEC, RSTC, SIGNEDA, SIGNEDB, SIGNEDC, RSTOUT, CEOUT, Z); //synthesis syn_black_box syn_lib_cell=1
    input [17:0] A;
    input [17:0] B;
    input [17:0] C;
    input CLK;
    input CEA;
    input RSTA;
    input CEB;
    input RSTB;
    input CEC;
    input RSTC;
    input SIGNEDA;
    input SIGNEDB;
    input SIGNEDC;
    input RSTOUT;
    input CEOUT;
    output [35:0] Z;
    parameter REGINPUTA = "REGISTER";
    parameter REGINPUTB = "REGISTER";
    parameter REGINPUTC = "REGISTER";
    parameter REGOUTPUT = "REGISTER";
    parameter GSR = "ENABLED";
    parameter RESETMODE = "SYNC";
endmodule

module MULTPREADD9X9(A, B, C, CLK, CEA, RSTA, CEB, RSTB, CEC, RSTC, SIGNEDA, SIGNEDB, SIGNEDC, RSTOUT, CEOUT, Z); //synthesis syn_black_box syn_lib_cell=1
    input [8:0] A;
    input [8:0] B;
    input [8:0] C;
    input CLK;
    input CEA;
    input RSTA;
    input CEB;
    input RSTB;
    input CEC;
    input RSTC;
    input SIGNEDA;
    input SIGNEDB;
    input SIGNEDC;
    input RSTOUT;
    input CEOUT;
    output [17:0] Z;
    parameter REGINPUTA = "REGISTER";
    parameter REGINPUTB = "REGISTER";
    parameter REGINPUTC = "REGISTER";
    parameter REGOUTPUT = "REGISTER";
    parameter GSR = "ENABLED";
    parameter RESETMODE = "SYNC";
endmodule

module ODDR71(D0, D1, D2, D3, D4, D5, D6, SCLK, RST, ECLK, Q); //synthesis syn_black_box syn_lib_cell=1
    input D0;
    input D1;
    input D2;
    input D3;
    input D4;
    input D5;
    input D6;
    input SCLK;
    input RST;
    input ECLK;
    output Q;
    parameter GSR = "ENABLED";
endmodule

module ODDRX1(D0, D1, SCLK, RST, Q); //synthesis syn_black_box syn_lib_cell=1
    input D0;
    input D1;
    input SCLK;
    input RST;
    output Q;
    parameter GSR = "ENABLED";
endmodule

module ODDRX2DQS(D0, D1, D2, D3, DQSW, ECLK, SCLK, RST, Q); //synthesis syn_black_box syn_lib_cell=1
    input D0;
    input D1;
    input D2;
    input D3;
    input DQSW;
    input ECLK;
    input SCLK;
    input RST;
    output Q;
    parameter GSR = "ENABLED";
endmodule

module ODDRX2DQ(D0, D1, D2, D3, DQSW270, ECLK, SCLK, RST, Q); //synthesis syn_black_box syn_lib_cell=1
    input D0;
    input D1;
    input D2;
    input D3;
    input DQSW270;
    input ECLK;
    input SCLK;
    input RST;
    output Q;
    parameter GSR = "ENABLED";
endmodule

module ODDRX2(D0, D1, D2, D3, SCLK, RST, ECLK, Q); //synthesis syn_black_box syn_lib_cell=1
    input D0;
    input D1;
    input D2;
    input D3;
    input SCLK;
    input RST;
    input ECLK;
    output Q;
    parameter GSR = "ENABLED";
endmodule

module ODDRX4DQS(D0, D1, D2, D3, D4, D5, D6, D7, DQSW, ECLK, SCLK, RST, Q); //synthesis syn_black_box syn_lib_cell=1
    input D0;
    input D1;
    input D2;
    input D3;
    input D4;
    input D5;
    input D6;
    input D7;
    input DQSW;
    input ECLK;
    input SCLK;
    input RST;
    output Q;
    parameter GSR = "ENABLED";
endmodule

module ODDRX4DQ(D0, D1, D2, D3, D4, D5, D6, D7, DQSW270, ECLK, SCLK, RST, Q); //synthesis syn_black_box syn_lib_cell=1
    input D0;
    input D1;
    input D2;
    input D3;
    input D4;
    input D5;
    input D6;
    input D7;
    input DQSW270;
    input ECLK;
    input SCLK;
    input RST;
    output Q;
    parameter GSR = "ENABLED";
endmodule

module ODDRX4(D0, D1, D2, D3, D4, D5, D6, D7, SCLK, RST, ECLK, Q); //synthesis syn_black_box syn_lib_cell=1
    input D0;
    input D1;
    input D2;
    input D3;
    input D4;
    input D5;
    input D6;
    input D7;
    input SCLK;
    input RST;
    input ECLK;
    output Q;
    parameter GSR = "ENABLED";
endmodule

module ODDRX5(D0, D1, D2, D3, D4, D5, D6, D7, D8, D9, SCLK, RST, ECLK, Q); //synthesis syn_black_box syn_lib_cell=1
    input D0;
    input D1;
    input D2;
    input D3;
    input D4;
    input D5;
    input D6;
    input D7;
    input D8;
    input D9;
    input SCLK;
    input RST;
    input ECLK;
    output Q;
    parameter GSR = "ENABLED";
endmodule

module OFD1P3BX(D, SP, CK, PD, Q); //synthesis syn_black_box syn_lib_cell=1
    input D;
    input SP;
    input CK;
    input PD;
    output Q;
    parameter GSR = "ENABLED";
endmodule

module OFD1P3DX(D, SP, CK, CD, Q); //synthesis syn_black_box syn_lib_cell=1
    input D;
    input SP;
    input CK;
    input CD;
    output Q;
    parameter GSR = "ENABLED";
endmodule

module OFD1P3IX(D, SP, CK, CD, Q); //synthesis syn_black_box syn_lib_cell=1
    input D;
    input SP;
    input CK;
    input CD;
    output Q;
    parameter GSR = "ENABLED";
endmodule

module OFD1P3JX(D, SP, CK, PD, Q); //synthesis syn_black_box syn_lib_cell=1
    input D;
    input SP;
    input CK;
    input PD;
    output Q;
    parameter GSR = "ENABLED";
endmodule

module OSHX2(D0, D1, ECLK, SCLK, RST, Q); //synthesis syn_black_box syn_lib_cell=1
    input D0;
    input D1;
    input ECLK;
    input SCLK;
    input RST;
    output Q;
    parameter GSR = "ENABLED";
endmodule

module OSHX4(D0, D1, D2, D3, ECLK, SCLK, RST, Q); //synthesis syn_black_box syn_lib_cell=1
    input D0;
    input D1;
    input D2;
    input D3;
    input ECLK;
    input SCLK;
    input RST;
    output Q;
    parameter GSR = "ENABLED";
endmodule

module PCIE(LMMICLK, LMMIRESET_N, LMMIREQUEST, LMMIWRRD_N, LMMIOFFSET, LMMIWDATA, LMMIRDATA, LMMIRDATAVALID, LMMIREADY, ACJNOUT, ACJPOUT, AUXCK, CKUSRI, CKUSRO, ECKIN, ECKIND2, ECKINDO, ERSTN, ERSTND2, ERXCKD2, ERXCKDO, ERXRSND2, ETXCKD2, ETXCKDO, ETXRSND2, FLR, FLRACK, MINTLEG, MINTO, PERSTN, PMCTRL, PMCTRLEN, PMDPAST, PRMSGSD, PRNOSNP, PRNSNPRE, PRSNOOP, PRSNPRE, PPBDREG, PPBDSEL, REXTCK, REXTRST, RSTUSRN, UDLLKUP, ULTSDIS, UPLLKUP, UTLLKUP, UCFGADDR, UCFGF, UCFGRDD, UCFGRDE, UCFGRDY, UCFGSERD, UCFGVD, UCFGWRBE, UCFGWRD, UCFGWRDN, USERAUPD, USERTRS, VRXCMDD, VRXCINIT, VRXCNH, VRXCNINF, VRXCRRE, VRXD, VRXDP, VRXEOP, VRXERR, VRXF, VRXRDY, VRXSEL, VRXSOP, VRXVD, VXCDINIT, VXCDNH, VTXCRRE, VXD, VXDP, VXEOP, VXEOPN, VXRDY, VXSOP, VXVD, TESTOUT, S0REFCKN, S0REFCKP, S0REFRET, S0REXT, S0RXN, S0RXP, S0TXN, S0TXP, CLKREQI, CLKREQO, CLKREQOE); //synthesis black_box_pad_pin="S0REFCKN,S0REFCKP,S0REFRET,S0REXT,S0RXN,S0RXP,S0TXN,S0TXP" syn_lib_cell=1
    input LMMICLK;
    input LMMIRESET_N;
    input LMMIREQUEST;
    input LMMIWRRD_N;
    input [14:0] LMMIOFFSET;
    input [31:0] LMMIWDATA;
    output [31:0] LMMIRDATA;
    output LMMIRDATAVALID;
    output LMMIREADY;
    output ACJNOUT;
    output ACJPOUT;
    input AUXCK;
    input CKUSRI;
    output CKUSRO;
    input ECKIN;
    input ECKIND2;
    output ECKINDO;
    input ERSTN;
    input ERSTND2;
    input ERXCKD2;
    output ERXCKDO;
    input ERXRSND2;
    input ETXCKD2;
    output ETXCKDO;
    input ETXRSND2;
    output [3:0] FLR;
    input [3:0] FLRACK;
    input [3:0] MINTLEG;
    output MINTO;
    input PERSTN;
    output [4:0] PMCTRL;
    output PMCTRLEN;
    input [4:0] PMDPAST;
    input PRMSGSD;
    input [12:0] PRNOSNP;
    input PRNSNPRE;
    input [12:0] PRSNOOP;
    input PRSNPRE;
    input [31:0] PPBDREG;
    output [7:0] PPBDSEL;
    input REXTCK;
    input REXTRST;
    input RSTUSRN;
    output UDLLKUP;
    input ULTSDIS;
    output UPLLKUP;
    output UTLLKUP;
    input [9:0] UCFGADDR;
    input [2:0] UCFGF;
    output [31:0] UCFGRDD;
    output UCFGRDE;
    output UCFGRDY;
    input UCFGSERD;
    input UCFGVD;
    input [3:0] UCFGWRBE;
    input [31:0] UCFGWRD;
    input UCFGWRDN;
    input USERAUPD;
    input [3:0] USERTRS;
    output [12:0] VRXCMDD;
    input VRXCINIT;
    input [11:0] VRXCNH;
    input VRXCNINF;
    input VRXCRRE;
    output [31:0] VRXD;
    output [3:0] VRXDP;
    output VRXEOP;
    output VRXERR;
    output [1:0] VRXF;
    input VRXRDY;
    output [1:0] VRXSEL;
    output VRXSOP;
    output VRXVD;
    output VXCDINIT;
    output [11:0] VXCDNH;
    output VTXCRRE;
    input [31:0] VXD;
    input [3:0] VXDP;
    input VXEOP;
    input VXEOPN;
    output VXRDY;
    input VXSOP;
    input VXVD;
    output [7:0] TESTOUT;
    input S0REFCKN;
    input S0REFCKP;
    input S0REFRET;
    input S0REXT;
    input S0RXN;
    input S0RXP;
    output S0TXN;
    output S0TXP;
    input CLKREQI;
    output CLKREQO;
    output CLKREQOE;
    parameter ENABLE_USER_CFG = "DISABLED";
    parameter PWDN_N = "DISABLED";
    parameter GSR = "ENABLED";
    parameter IDDQ_PCS = "DISABLED";
    parameter PHY_MODE = "0b0000";
    parameter ALT_CLK_SEL_VCC = "PAD";
    parameter L0S_ADJ = "0b00000110000000";
    parameter L0S_EXIT_LATENCY = "MORE_4_US";
    parameter L1_EXIT_LATENCY = "MORE_64_US";
    parameter CALIB_3DB = "ENABLED";
    parameter DB_UPSTREAM = "6DB";
    parameter ERR_REC_ENTRY_SEL = "RCVRY_AFTER";
    parameter A_CHNGD_MAX = "0b100";
    parameter A0_FORCE = "DISABLED";
    parameter A0_FREEZE = "DISABLED";
    parameter A0_INIT = "0b000000";
    parameter A0DIR_VAL = "DISABLED";
    parameter A1_FORCE = "DISABLED";
    parameter A1_FREEZE = "DISABLED";
    parameter A1_INIT = "0b000000";
    parameter A1DIR_VAL = "DISABLED";
    parameter A2_FORCE = "DISABLED";
    parameter A2_FREEZE = "DISABLED";
    parameter A2_INIT = "0b000000";
    parameter A2GAIN_CALIB = "0b100110";
    parameter ACJTAG_REG = "0b00";
    parameter ADDR_LIMIT_PRE_MTHD_CTRL = "0b0100";
    parameter ADDR_LIMIT_TABLE_MTHD_CTRL = "0b00101";
    parameter ADIR_OVR = "DISABLED";
    parameter ADV_CH_CD_SEL = "IMPLEMENT_CH";
    parameter ADV_TARGET_LINK_SPEED_USPORT_A = "DISABLED";
    parameter ADV_TARGET_LINK_SPEED_USPORT_B = "DISABLED";
    parameter ADV_TARGET_LINK_SPEED_USPORT_C = "DISABLED";
    parameter ADV_TARGET_LINK_SPEED_USPORT_D = "DISABLED";
    parameter ADVANCE = "DISABLED";
    parameter ALERT_ENABLE = "0b000";
    parameter ALMOST_EMPTY_10B = "0b001110";
    parameter MID_VALUE_10B = "0b011110";
    parameter ALMOST_EMPTY_20B = "0b001111";
    parameter ALMOST_EMPTY_GEN3 = "0b001100";
    parameter ALMOST_FULL_10B = "0b110000";
    parameter ALMOST_FULL_20B = "0b011000";
    parameter ALMOST_FULL_GEN3 = "0b010110";
    parameter ARRAY_DA = "0b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter ARRAY_MT = "0b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000011100000000000010000000000000001001000000000000011000000000000001010000000000000100";
    parameter ARXCDRICP_RATE0 = "0b011";
    parameter ARXCDRICP_RATE1 = "0b011";
    parameter ARXCDRICP_RATE2 = "0b011";
    parameter ARXDMPWRDWN = "DISABLED";
    parameter ARXDPPWRDN = "DISABLED";
    parameter ARXEOM_PWRDN = "POWERED_DOWN";
    parameter ARXICP_RATE0 = "0b011";
    parameter ARXICP_RATE1 = "0b011";
    parameter ARXICP_RATE2 = "0b011";
    parameter ARXOVR_OUT = "DISABLED";
    parameter ARXRSACTAT = "0b0001";
    parameter ARXRSAPTAT = "0b1000";
    parameter ARXRSVCTL = "0b00000000";
    parameter ARXSEL_OUT = "DISABLED";
    parameter ASPM_L1_1_SUPPORTED = "SUPPORTED";
    parameter ASPM_L1_2_SUPPORTED = "SUPPORTED";
    parameter ASPM_SUPPORT = "L0S_AND_L1_SUPPORTED";
    parameter ATTENTION_BUTTON_PRESENT = "NOT_SUPPORTED";
    parameter ATTENTION_INDICATOR_PRESENT = "NOT_SUPPORTED";
    parameter ATXICP_RATE0 = "0b101";
    parameter ATXICP_RATE1 = "0b101";
    parameter AUTO_SHIFT = "ENABLED";
    parameter AUX_CURRENT = "SELF_POWERED";
    parameter AUXCLK1US_MAX = "0b00001001";
    parameter AUXIDL_MAX = "0b00000100";
    parameter BAR_INDEX_CFG0_A = "0b000";
    parameter BAR_INDEX_CFG0_B = "0b000";
    parameter BAR_INDEX_CFG0_C = "0b000";
    parameter BAR_INDEX_CFG0_D = "0b000";
    parameter BAR_INDEX_CFG1_A = "0b001";
    parameter BAR_INDEX_CFG1_B = "0b001";
    parameter BAR_INDEX_CFG1_C = "0b001";
    parameter BAR_INDEX_CFG1_D = "0b001";
    parameter BAR_INDEX_CFG2_A = "0b010";
    parameter BAR_INDEX_CFG2_B = "0b010";
    parameter BAR_INDEX_CFG2_C = "0b010";
    parameter BAR_INDEX_CFG2_D = "0b010";
    parameter BAR_INDEX_CFG3_A = "0b011";
    parameter BAR_INDEX_CFG3_B = "0b011";
    parameter BAR_INDEX_CFG3_C = "0b011";
    parameter BAR_INDEX_CFG3_D = "0b011";
    parameter BAR_INDEX_CFG4_A = "0b100";
    parameter BAR_INDEX_CFG4_B = "0b100";
    parameter BAR_INDEX_CFG4_C = "0b100";
    parameter BAR_INDEX_CFG4_D = "0b100";
    parameter BAR_INDEX_CFG5_A = "0b101";
    parameter BAR_INDEX_CFG5_B = "0b101";
    parameter BAR_INDEX_CFG5_C = "0b101";
    parameter BAR_INDEX_CFG5_D = "0b101";
    parameter BIR_MSIX_PBA_A = "BAR0";
    parameter BIR_MSIX_PBA_B = "BAR0";
    parameter BIR_MSIX_PBA_C = "BAR0";
    parameter BIR_MSIX_PBA_D = "BAR0";
    parameter BIR_MSIX_TABLE_A = "BAR0";
    parameter BIR_MSIX_TABLE_B = "BAR0";
    parameter BIR_MSIX_TABLE_C = "BAR0";
    parameter BIR_MSIX_TABLE_D = "BAR0";
    parameter BYP_AVG = "USED";
    parameter BYPASS = "PERFORM_RECEIVER_DETECTION";
    parameter BYPASS_ADDR_DEC = "NORMAL";
    parameter CALIB_SETTLE_MAX = "0b001";
    parameter CALIB_STABLE_MAX = "0b11000";
    parameter CAPABILITY_VERSION = "0b0010";
    parameter CDR_ERR = "DISABLED";
    parameter CDR_P1 = "CDR_PLL_RESET";
    parameter CDR_PLL_DELTA = "0P4_PERCENT";
    parameter CDR_REFERENCE = "0b00";
    parameter CDRPLL_CMP_MAX = "0b00010100";
    parameter CDRPLL_CNT_MAX = "0b00000100";
    parameter CDRPLL_PRE_RXEQ_COARSE_TIMER = "0b01010000";
    parameter CDRPLL_PRE_RXEQ_FINE_TIMER = "0b10110100";
    parameter CDRPLL_PST_RXEQ_COARSE_TIMER = "0b01000000";
    parameter CDRPLL_PST_RXEQ_FINE_TIMER = "0b01000010";
    parameter CFG_A_BAR0 = "0b11111111111111110000000000001100";
    parameter CFG_A_BAR1 = "0b11111111111111111111111111111111";
    parameter CFG_A_BAR2 = "0b11111111111111111110000000001100";
    parameter CFG_A_BAR3 = "0b11111111111111111111111111111111";
    parameter CFG_A_BAR4 = "0b11111111111111111110000000001100";
    parameter CFG_A_BAR5 = "0b11111111111111111111111111111111";
    parameter CFG_B_BAR0 = "0b11111111111111110000000000001100";
    parameter CFG_B_BAR1 = "0b11111111111111111111111111111111";
    parameter CFG_B_BAR2 = "0b11111111111111111110000000001100";
    parameter CFG_B_BAR3 = "0b11111111111111111111111111111111";
    parameter CFG_B_BAR4 = "0b11111111111111111110000000001100";
    parameter CFG_B_BAR5 = "0b11111111111111111111111111111111";
    parameter CFG_C_BAR0 = "0b11111111111111110000000000001100";
    parameter CFG_C_BAR1 = "0b11111111111111111111111111111111";
    parameter CFG_C_BAR2 = "0b11111111111111111110000000001100";
    parameter CFG_C_BAR3 = "0b11111111111111111111111111111111";
    parameter CFG_C_BAR4 = "0b11111111111111111110000000001100";
    parameter CFG_C_BAR5 = "0b11111111111111111111111111111111";
    parameter CFG_D_BAR0 = "0b11111111111111110000000000001100";
    parameter CFG_D_BAR1 = "0b11111111111111111111111111111111";
    parameter CFG_D_BAR2 = "0b11111111111111111110000000001100";
    parameter CFG_D_BAR3 = "0b11111111111111111111111111111111";
    parameter CFG_D_BAR4 = "0b11111111111111111110000000001100";
    parameter CFG_D_BAR5 = "0b11111111111111111111111111111111";
    parameter CFG_EXP_ROM_A = "0b00000000000000000000000000000000";
    parameter CFG_EXP_ROM_B = "0b00000000000000000000000000000000";
    parameter CFG_EXP_ROM_C = "0b00000000000000000000000000000000";
    parameter CFG_EXP_ROM_D = "0b00000000000000000000000000000000";
    parameter CIS_POINTER_CARDBUS_A = "0b00000000000000000000000000000000";
    parameter CIS_POINTER_CARDBUS_B = "0b00000000000000000000000000000000";
    parameter CIS_POINTER_CARDBUS_C = "0b00000000000000000000000000000000";
    parameter CIS_POINTER_CARDBUS_D = "0b00000000000000000000000000000000";
    parameter CLASS_CODE_ID3A = "0b000100011000000000000000";
    parameter CLASS_CODE_ID3B = "0b000100011000000000000000";
    parameter CLASS_CODE_ID3C = "0b000100011000000000000000";
    parameter CLASS_CODE_ID3D = "0b000100011000000000000000";
    parameter CM_RESTORE_TIME = "0b00000000";
    parameter CNT250NS_MAX = "0b001111100";
    parameter COARSE_GAIN = "DISABLED";
    parameter COEF_EN_LPBK_MASTER = "OTHERWISE";
    parameter COEF_EN_LPBK_SLAVE = "OTHERWISE";
    parameter COEF_ENABLE = "DETERMINE_LOCAL_PHY";
    parameter COEF_EQTX_FORCE = "0b000000000000000000";
    parameter COEF_LPBK_MASTER = "0b000000000000000000";
    parameter COEF_LPBK_SLAVE = "0b000000000000000000";
    parameter COEF0_POST = "0b000101";
    parameter COEF0_POST_CURSOR = "0b000000";
    parameter COEF0_PRE = "0b000000";
    parameter COEF0_PRE_CURSOR = "0b000000";
    parameter COEF1_POST = "0b000011";
    parameter COEF1_POST_CURSOR = "0b000000";
    parameter COEF1_PRE = "0b000000";
    parameter COEF1_PRE_CURSOR = "0b000000";
    parameter COEF10_POST = "0b000111";
    parameter COEF10_PRE = "0b000000";
    parameter COEF2_POST = "0b000100";
    parameter COEF2_POST_CURSOR = "0b000000";
    parameter COEF2_PRE = "0b000000";
    parameter COEF2_PRE_CURSOR = "0b000000";
    parameter COEF3_POST = "0b000010";
    parameter COEF3_POST_CURSOR = "0b000000";
    parameter COEF3_PRE = "0b000000";
    parameter COEF3_PRE_CURSOR = "0b000000";
    parameter COEF4_POST = "0b000000";
    parameter COEF4_PRE = "0b000000";
    parameter COEF5_POST = "0b000000";
    parameter COEF5_PRE = "0b000001";
    parameter COEF6_POST = "0b000000";
    parameter COEF6_PRE = "0b000010";
    parameter COEF7_POST = "0b000100";
    parameter COEF7_PRE = "0b000011";
    parameter COEF8_POST = "0b000011";
    parameter COEF8_PRE = "0b000010";
    parameter COEF9_POST = "0b000000";
    parameter COEF9_PRE = "0b000011";
    parameter COMP_128_SUPPORTED = "ENABLED";
    parameter COMP_32_SUPPORTED = "ENABLED";
    parameter COMP_64_SUPPORTED = "ENABLED";
    parameter COMPLETE = "DISABLED";
    parameter CONV_METHOD = "COMPUTE_PCIE_SPEC";
    parameter CORE_BYPASS = "NORMAL";
    parameter CORE_EN = "ENABLED";
    parameter COUNT_ACK_TO_NAK = "0b00000000";
    parameter CPL_TIMEOUT_DISABLE_SUPPORTED = "SUPPORTED";
    parameter CPL_TIMEOUT_RANGES_SUPPORTED = "NOT_SUPPORTED";
    parameter CRS_ENABLE = "DISABLED";
    parameter CSTAT_DATA_SCALE = "UNKNOWN_SCALE";
    parameter CSTAT_DATA_SELECT = "D0_POWER_CONSUMED";
    parameter CTLE_SETTLE = "0b100";
    parameter CTLEBIAS_1 = "0b1000";
    parameter ATXICP_RATE2 = "0b100";
    parameter CTLEBYPASS = "DISABLED";
    parameter CUR_FOM = "NUMBER_OF_CLOCK";
    parameter CUR_FOM_AVG = "0b101";
    parameter CUST_AUTO = "DISABLED";
    parameter CUST_CHK = "SET";
    parameter CUST_SEL = "DISABLED";
    parameter CUST_SKIP = "DISABLED";
    parameter CUST_TYP = "0b000";
    parameter CUSTOM_PATTERN = "0b00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter D1_SUPPORT = "SUPPORTED";
    parameter D2_SUPPORT = "SUPPORTED";
    parameter DATA_INJECT = "0b00000000000000000000000000000000";
    parameter DATA_PM = "0b00000000";
    parameter DEEMPH_5G_3_5DB_6DB_N = "6DB";
    parameter DEEMPH_5G_ENABLE = "DISABLED";
    parameter DEEMPH_LPBK_MASTER = "6P0DB";
    parameter DEEMPH_LPBK_SLAVE = "6P0DB";
    parameter DEVICE_ID_ID1A = "0b1110000000000100";
    parameter DEVICE_ID_ID1B = "0b1110000000000100";
    parameter DEVICE_ID_ID1C = "0b1110000000000100";
    parameter DEVICE_ID_ID1D = "0b1110000000000100";
    parameter DEVICE_PORT_TYPE = "PCIE_ENDPOINT";
    parameter DFE_BIAS = "0b0001";
    parameter DFE_PWDN = "DISABLED";
    parameter DIR_PRE_GAIN = "0b00";
    parameter DIR_PST_GAIN = "0b01";
    parameter DIS_ARI_CAP = "ENABLED";
    parameter DIS_CSR_RST = "DISABLED";
    parameter DIS_INTERRUPT = "ENABLED";
    parameter DIS_INTERRUPT_B = "ENABLED";
    parameter DIS_INTERRUPT_C = "ENABLED";
    parameter DIS_INTERRUPT_D = "ENABLED";
    parameter DIS_MSI_CAP = "ENABLED";
    parameter DIS_MSI_CAP_B = "ENABLED";
    parameter DIS_MSI_CAP_C = "ENABLED";
    parameter DIS_MSI_CAP_D = "ENABLED";
    parameter DIS_MSIX_CAP = "ENABLED";
    parameter DIS_MSIX_CAP_B = "ENABLED";
    parameter DIS_MSIX_CAP_C = "ENABLED";
    parameter DIS_MSIX_CAP_D = "ENABLED";
    parameter DISABLE_FLR_CAPABILITY = "ENABLED";
    parameter DLLP_CRC_ERR_ENABLE = "DISABLED";
    parameter DLLP_CRC_ERR_RATE = "0b000000000000";
    parameter DLLP_INJECT_ENABLE = "DISABLED";
    parameter DOUBLE_TX_DATA_VALID = "ONE_CLK_EVERY_64_CLKS";
    parameter DOWNSTREAM_EQ_SKIP_PHASE_2_3 = "NORMAL_OPERATION";
    parameter DS_DRIVE_CLKREQ = "ENABLED";
    parameter DS_PORT_RX_PRESET_HINT = "0b001";
    parameter DS_PORT_TX_PRESET = "0b0011";
    parameter DS_US_N_PORTTYPE = "UPSTREAM";
    parameter DSI = "NO_DSI_NECESSARY";
    parameter DSP_DIR = "ANALYSIS_OF_DATA_BY_DSP";
    parameter DSPDIR_PRESGN = "0b11110000";
    parameter DSPDIR_PREVAL = "0b00011000";
    parameter DSPDIR_PSTSGN0 = "0b11111111";
    parameter DSPDIR_PSTSGN1 = "0b00000000";
    parameter DSPDIR_PSTVAL0 = "0b00000010";
    parameter DSPDIR_PSTVAL1 = "0b01000000";
    parameter EARLY_RX_EVAL = "RX_SIGNAL_AFTER_TS1";
    parameter ECRC_GEN_CHK_CAPABLE = "SUPPORTED";
    parameter EFF_LPBK = "PASSED";
    parameter EI4 = "EI_IV";
    parameter EM_INTERLOCK_PRESENT = "NOT_SUPPORTED";
    parameter EN = "DISABLED";
    parameter EN_ACK_TO_DIV = "ACK_SPEC";
    parameter EN_ACK_TO_NAK = "DO_NOTHING";
    parameter EN_ACS_VIOLATION = "DISABLED";
    parameter EN_ASPM_L0S = "ENABLED";
    parameter EN_ASPM_L1 = "ENABLED";
    parameter EN_ATOMIC_OP_CAP = "ENABLED";
    parameter EN_ATOMICOP_EGRESS_BLOCKED = "DISABLED";
    parameter EN_ATS_CAP = "ENABLED";
    parameter EN_BDGT_CAP = "DISABLED";
    parameter EN_CAP = "ENABLED";
    parameter EN_CAP_B = "ENABLED";
    parameter EN_CAP_C = "ENABLED";
    parameter EN_CAP_D = "ENABLED";
    parameter EN_COMPLETER_ABORT = "DISABLED";
    parameter EN_COMPLETION_TIMEOUT = "ENABLED";
    parameter EN_CORR_INTERNAL_ERROR = "DISABLED";
    parameter EN_DPA_CAP = "DISABLED";
    parameter EN_DRCT_SCR_OFF = "OTHERWISE";
    parameter EN_DRCT_TO_LPBK = "OTHERWISE";
    parameter EN_EQTX_OVERRIDE = "PIPE_LOCAL_FS_AND_PIPE_LOCAL_LF";
    parameter EN_FORCE_SCR_OFF_FAST = "OTHERWISE";
    parameter EN_L1 = "ENABLED";
    parameter EN_L1PMSS_CAP = "ENABLED";
    parameter EN_L2 = "ENABLED";
    parameter EN_LPBK_ERR_RST = "MASTER_LPBK_INCREMENT";
    parameter EN_LTR_CAP = "ENABLED";
    parameter EN_MC_BLOCKED_TLP = "DISABLED";
    parameter EN_NWL_VSEC_CAP = "ENABLED";
    parameter EN_PORT_DIS = "DISABLED";
    parameter EN_PORT_INTLEG = "ENABLED";
    parameter EN_RBAR_CAP_A = "ENABLED";
    parameter EN_RBAR_CAP_B = "ENABLED";
    parameter EN_RBAR_CAP_C = "ENABLED";
    parameter EN_RBAR_CAP_D = "ENABLED";
    parameter EN_RECEIVER_OVERFLOW = "DISABLED";
    parameter EN_SELF_XLINK = "OTHERWISE";
    parameter EN_SURPRISE_DOWN_ERROR = "DISABLED";
    parameter EN_TLP_PREFIX_BLOCKED = "DISABLED";
    parameter EN_UCORR_INTERNAL_ERROR = "DISABLED";
    parameter EN_USER_WRITE = "READ_WRITE_ACCESS";
    parameter END_END_PREFIXES_SUPPORTED = "NOT_SUPPORTED";
    parameter END_ON_HOLD = "YES_EXIT_ON_HOLD";
    parameter ENDCALIB_MAX = "0b10000100";
    parameter ENDPOINT_L0S_ACCEPTABLE_LATENCY = "MAX_64_NS";
    parameter ENDPOINT_L1_ACCEPTABLE_LATENCY = "MAX_1_US";
    parameter ENTRY_TIME_ASPM_L0S = "0b0000000000000000";
    parameter ENTRY_TIME_ASPM_L1 = "0b0000000000000000";
    parameter EOM_TIME = "0b0000000000000000";
    parameter EOM0DIR = "SELECT_DIR_1";
    parameter EOM1DIR = "SELECT_DIR_0";
    parameter EOMCTRL0_LOW = "DISABLED";
    parameter EOMDIVDIS = "DISABLED";
    parameter EOMMODE = "0b00";
    parameter EOMRDSEL = "DISABLED";
    parameter EOMSTART = "DISABLED";
    parameter EOMX = "0b000000";
    parameter EOMX_UPDATE_CNT_VALUE = "0b0011111";
    parameter EOMY = "0b00000000";
    parameter ERRCNT_DEC = "0b00100000";
    parameter ERRCNT_THR = "0b1000";
    parameter ES_PWDN = "DISABLED";
    parameter EVAL_RST = "DISABLED";
    parameter EXCLUDE_L0 = "INCLUDE";
    parameter EXCLUDE_CFG_COMPLETE = "INCLUDE";
    parameter EXCLUDE_CFG_IDLE = "INCLUDE";
    parameter EXCLUDE_LOOPBACK_MASTER = "INCLUDE";
    parameter EXCLUDE_REC_IDLE = "INCLUDE";
    parameter EXCLUDE_REC_RCVR_CFG = "INCLUDE";
    parameter EXIT_DIRECT_TO_DETECT = "DO_NOT_EXIT_TO_DETECT";
    parameter EXT_CONTROL = "DISABLED";
    parameter EXTENDED_TAG_FIELD_EN_DEFAULT = "EIGHT_BIT";
    parameter EXTENDED_TAG_FIELD_SUPPORTED = "EIGHT_BIT";
    parameter F_ARXCTLEDIR = "IGNORED";
    parameter F_ARXCTLENULL = "0b0000";
    parameter F_ARXDMDIR = "DISABLED";
    parameter F_ARXDMNULL = "0b00000";
    parameter F_ARXEOMDIR = "IGNORED";
    parameter F_ARXEOMNULL = "0b00000";
    parameter F_ARXESDIR = "IGNORED";
    parameter F_ARXESNULL = "0b00000";
    parameter F_ARXTDIR = "IGNORED";
    parameter F_ARXTNULL = "0b00000";
    parameter F_ASCHCAL = "IGNORED";
    parameter F_ASCHDIR = "IGNORED";
    parameter F_ASCHNULL = "0b0000";
    parameter FAIL_LIMIT_ERR = "RXEQ_NOT_FAIL";
    parameter FAST = "L0";
    parameter FC_UPDATE_TIMER_DISABLE = "ENABLED";
    parameter FC_UPDATE_TIMER_DIV = "PCIE_REC_VALUES";
    parameter FILTER = "0b1001";
    parameter FINE_GAIN = "DISABLED";
    parameter FOM_COMPARE = "0b00000000";
    parameter FOM_HIRES = "DISABLED";
    parameter FOM_ITERCNT = "0b101";
    parameter FOM_THR = "0b0100";
    parameter FORCE_ATXDRA = "0b000000000000000000000";
    parameter FORCE_ATXDRP = "0b000000000000000000000";
    parameter FORCE_ATXDRR = "0b000000000000000000000";
    parameter FORCE_ATXDRT = "0b000000000000000000000";
    parameter FORCE_DIR_RSLT = "0b000000";
    parameter FORCE_FOM_RSLT = "0b00000000";
    parameter FORCE_IDLE = "DISABLED";
    parameter FORCE_RX_DETECT = "DISABLED";
    parameter FORCE_SIGNAL = "DISABLED";
    parameter FREQ_LOCK = "DISABLED";
    parameter FS = "0b110000";
    parameter GAIN_TIMER1 = "0b0101";
    parameter GEN12_ENA_POST_A0 = "DISABLED";
    parameter GEN12_ENA_POST_A1A2 = "DISABLED";
    parameter GEN12_ENA_PREA0 = "DISABLED";
    parameter GEN3_ENA_POST_A0 = "ENABLED";
    parameter GEN3_ENA_POST_A1A2 = "ENABLED";
    parameter GEN3_ENA_PREA0 = "ENABLED";
    parameter GLOBAL_INVAL_SUPPORT = "ENABLED";
    parameter HINT = "0b000";
    parameter HINT0_3DB = "ENABLED";
    parameter HINT0_A0GAIN = "0b111";
    parameter HINT0_A2GAIN = "0b111";
    parameter HINT1_3DB = "ENABLED";
    parameter HINT1_A0GAIN = "0b011";
    parameter HINT1_A2GAIN = "0b101";
    parameter HINT2_3DB = "ENABLED";
    parameter HINT2_A0GAIN = "0b011";
    parameter HINT2_A2GAIN = "0b111";
    parameter HINT3_3DB = "ENABLED";
    parameter HINT3_A0GAIN = "0b000";
    parameter HINT3_A2GAIN = "0b111";
    parameter HINT4_3DB = "DISABLED";
    parameter HINT4_A0GAIN = "0b111";
    parameter HINT4_A2GAIN = "0b111";
    parameter HINT5_3DB = "DISABLED";
    parameter HINT5_A0GAIN = "0b011";
    parameter HINT5_A2GAIN = "0b101";
    parameter HINT6_3DB = "DISABLED";
    parameter HINT6_A0GAIN = "0b011";
    parameter HINT6_A2GAIN = "0b111";
    parameter HINT7_3DB = "DISABLED";
    parameter HINT7_A0GAIN = "0b000";
    parameter HINT7_A2GAIN = "0b111";
    parameter HINT7_OVR = "DISABLED";
    parameter HLD_RST = "WRITE_1";
    parameter HOT_PLUG_CAPABLE = "NOT_SUPPORTED";
    parameter HOT_PLUG_SURPRISE = "NOT_POSSIBLE";
    parameter ID_DS_PORT = "0b0000000000000000";
    parameter ID_NWL_VSEC_CAP = "0b0000000000000001";
    parameter IGNORE_ECRC = "DISABLED";
    parameter IGNORE_POISON = "ENABLED";
    parameter INDICATOR = "0b00000000000000000000000000000000";
    parameter INHIBIT = "PERFORM_RECEIVER_DETECTION";
    parameter INJECT_DATA_ERROR_0 = "DISABLED";
    parameter INJECT_DATA_ERROR_1 = "DISABLED";
    parameter INJECT_DATA_ERROR_2 = "DISABLED";
    parameter INJECT_DATA_ERROR_3 = "DISABLED";
    parameter INJECT_DATA_ERROR_EN = "DISABLED";
    parameter INJECT_ERR_LANE_SELECT_0 = "DISABLED";
    parameter INJECT_ERR_LANE_SELECT_1 = "DISABLED";
    parameter INJECT_ERR_LANE_SELECT_2 = "DISABLED";
    parameter INJECT_ERR_LANE_SELECT_3 = "DISABLED";
    parameter INJECT_RX_1BIT_DATA_ERR = "DISABLED";
    parameter INJECT_RX_2BIT_DATA_ERR = "DISABLED";
    parameter INJECT_RX_SKP_ERR = "DISABLED";
    parameter INJECT_RX_VALID_ERR = "DISABLED";
    parameter INT_CLR = "DISABLED";
    parameter INT_EN = "DISABLED";
    parameter INTERRUPT_MESSAGE_NUMBER = "0b00000";
    parameter INVAL_Q_DEPTH = "0b00000";
    parameter ITERATION_MAX = "0b000000";
    parameter L1_ENTER_PLL_RESET_TIME = "0b100";
    parameter L1_EXIT_PLL_LOCK_TIME = "0b01110";
    parameter L1PM_SUPPORTED = "SUPPORTED";
    parameter L2_D3HOT_ENABLE = "DISABLED";
    parameter LANE_SELECT = "0b0000";
    parameter LF = "0b001000";
    parameter LF_PHY = "0b001010";
    parameter LINK_LANE = "ENABLED";
    parameter LPBK_EN = "DISABLED";
    parameter LW_START_UPDN_ACK_EN = "DISABLED";
    parameter LW_START_UPDN_COUNT = "0b000011111010";
    parameter LW_START_UPDN_EIE_EN = "DISABLED";
    parameter LW_START_UPDN_EN_DIR_DS = "DO_NOT_ASSERT";
    parameter LW_START_UPDN_END_DELAY = "0b1001";
    parameter LW_START_UPDN_RATE_EN_16G = "DISABLED";
    parameter LW_START_UPDN_RATE_EN_2P5G = "ENABLED";
    parameter LW_START_UPDN_RATE_EN_5G = "ENABLED";
    parameter LW_START_UPDN_RATE_EN_8G = "ENABLED";
    parameter LW_START_UPDN_START_DELAY = "0b1000";
    parameter LW_START_UPDN_TIMER_EN = "DISABLED";
    parameter MARGIN_ENABLE = "PCIE_SPEC";
    parameter MARGIN_VALUE = "0b000";
    parameter MASK_0 = "SKIP_RCVR_DETECTION";
    parameter MASK_1 = "SKIP_RCVR_DETECTION";
    parameter MASK_2 = "SKIP_RCVR_DETECTION";
    parameter MASK_3 = "SKIP_RCVR_DETECTION";
    parameter MAX_LINK_WIDTH = "1_LANE";
    parameter MAX_SPEED = "8G";
    parameter MAX_VAR = "0b00100";
    parameter MERGE_LMMI_RDATA = "DISABLED";
    parameter METHOD_FMERIT_CTRL = "STEP_PCIE_TX_PRESETS";
    parameter METHOD_TX_CRED_CLEANUP = "HEADER";
    parameter MGMT_INTLEG = "0b0000";
    parameter MGMT_LTSSM_DIS = "DISABLED";
    parameter MID_VALUE_20B = "0b010100";
    parameter MID_VALUE_GEN3 = "0b001110";
    parameter MIN_SPEED = "2P5G";
    parameter MIN_TIME = "0_MS";
    parameter MIN_TIME_CFG = "4US";
    parameter MIX_DIR = "DISABLED";
    parameter MODE_BFF = "RESTART";
    parameter MRL_SENSOR_PRESENT = "NOT_SUPPORTED";
    parameter MULT_ENABLE = "RECOMMENDED_VALUES";
    parameter MULT_MESSAGE_CAPABLE_MSICAP_A = "EIGHT";
    parameter MULT_MESSAGE_CAPABLE_MSICAP_B = "EIGHT";
    parameter MULT_MESSAGE_CAPABLE_MSICAP_C = "EIGHT";
    parameter MULT_MESSAGE_CAPABLE_MSICAP_D = "EIGHT";
    parameter NFTS = "0b11111111";
    parameter NO_COMMAND_COMPLETED_SUPPORT = "SW_NOTIF_PROVIDED";
    parameter NO_FCMP = "DISABLED";
    parameter NO_REMOTE_CHANGE = "DISABLED";
    parameter NO_TX_IDLE_DELAY = "DATA_VALID_GAP";
    parameter NUM_LANES = "1_LANE";
    parameter NUMBER_DSLINK = "0b00000";
    parameter NUMHI_A = "0b00000000000000000000000000000000";
    parameter NUMHI_B = "0b00000000000000000000000000000000";
    parameter NUMHI_C = "0b00000000000000000000000000000000";
    parameter NUMHI_D = "0b00000000000000000000000000000000";
    parameter NUMHOLD = "SINGLE_HOLD_RESPONSE";
    parameter NUMLO_A = "0b00000000000000000000000000000000";
    parameter NUMLO_B = "0b00000000000000000000000000000000";
    parameter NUMLO_C = "0b00000000000000000000000000000000";
    parameter NUMLO_D = "0b00000000000000000000000000000000";
    parameter OBFF_SUPPORTED = "NOT_SUPPORTED";
    parameter OFFSET_MSIX_PBA_A = "0b00000000000000000111000000000";
    parameter OFFSET_MSIX_PBA_B = "0b00000000000000000111000000000";
    parameter OFFSET_MSIX_PBA_C = "0b00000000000000000111000000000";
    parameter OFFSET_MSIX_PBA_D = "0b00000000000000000111000000000";
    parameter OFFSET_MSIX_TABLE_A = "0b00000000000000000110000000000";
    parameter OFFSET_MSIX_TABLE_B = "0b00000000000000000110000000000";
    parameter OFFSET_MSIX_TABLE_C = "0b00000000000000000110000000000";
    parameter OFFSET_MSIX_TABLE_D = "0b00000000000000000110000000000";
    parameter OVER_CTLE = "DISABLED";
    parameter OVER_RX = "DISABLED";
    parameter OVER_RXDM = "DISABLED";
    parameter OVER_RXDP = "DISABLED";
    parameter OVER_RXES = "DISABLED";
    parameter OVER_RXT = "DISABLED";
    parameter OVER_SCH = "DISABLED";
    parameter OVER_TX = "DISABLED";
    parameter OVERRIDE = "DISABLED";
    parameter OVR_CDR = "DISABLED";
    parameter OVR_DIR = "DISABLED";
    parameter OVR_FOM = "DISABLED";
    parameter OVR_GAIN3DB = "ENABLED";
    parameter OVR_HINT3DB = "ENABLED";
    parameter P_CLK_PERIOD = "0b0000111110100000";
    parameter PAR_LPBK = "DISABLED";
    parameter PAS = "10X";
    parameter PATTERN_0 = "UNSCRAMBLED";
    parameter PATTERN_1 = "UNSCRAMBLED";
    parameter PATTERN_2 = "UNSCRAMBLED";
    parameter PCIPM_L1_1_SUPPORTED = "SUPPORTED";
    parameter PCIPM_L1_2_SUPPORTED = "SUPPORTED";
    parameter PERIOD_SRIS_128B130B = "0b000000";
    parameter PERIOD_SRIS_8B10B = "0b00000000";
    parameter PERIOD_SRNS_128B130B = "0b00000000";
    parameter PERIOD_SRNS_8B10B = "0b00000000";
    parameter PHANTOM_FUNCTIONS_SUPPORTED = "NO_FUNCTION_BITS";
    parameter PHYSICAL_SLOT_NUMBER = "0b0000000000001";
    parameter PIN_INTERRUPT_A = "INTA";
    parameter PIN_INTERRUPT_B = "INTA";
    parameter PIN_INTERRUPT_C = "INTA";
    parameter PIN_INTERRUPT_D = "INTA";
    parameter PIPE_TX_SWING = "FULL_SWING";
    parameter PLESIO_LPBK = "DISABLED";
    parameter PM_REDUCE_TIMEOUTS = "DISABLED";
    parameter PMA_DRIVEN_MODE = "PCS_DRIVEN";
    parameter PMCSR_B2_B3_SUPPORT = "DISABLED";
    parameter PMCSR_BUS_P_C_EN = "DISABLED";
    parameter PME_CLOCK = "DISABLED";
    parameter PME_SUPPORT = "0b11111";
    parameter PMFF_ALL = "DISABLED";
    parameter PORT_CM_RESTORE_TIME = "0b00000000";
    parameter PORT_NUMBER = "0b00000000";
    parameter PORT_TPOWER_ON_SCALE = "2_US";
    parameter PORT_TPOWER_ON_VALUE = "0b00000";
    parameter POST = "0b000000";
    parameter POST_A0COEF = "0b001";
    parameter POST_A1COEF = "0b001";
    parameter POST_A2COEF = "0b001";
    parameter POST_CURSOR_LIMIT = "0b100000";
    parameter POST_CURSOR_STEP_SIZE = "0b001000";
    parameter POST_ITERCNT = "0b100";
    parameter POST_STEP = "STEP_SIZE_4";
    parameter POWER_CONTROLLER_PRESENT = "NOT_SUPPORTED";
    parameter POWER_INDICATOR_PRESENT = "NOT_SUPPORTED";
    parameter POWER_REQUIRED = "AUX_POWER_NOT_REQUIRED";
    parameter PRBS_CHK = "DISABLED";
    parameter PRBS_GEN = "DISABLED";
    parameter PRBS_TYP = "PRBS7";
    parameter PRE = "0b000000";
    parameter PRE_A0COEF = "0b101";
    parameter PRE_A1COEF = "0b101";
    parameter PRE_A2COEF = "0b101";
    parameter PRE_CURSOR_LIMIT = "0b010000";
    parameter PRE_CURSOR_STEP_SIZE = "0b000100";
    parameter PRE_FOM = "ENABLED";
    parameter PRE_FOM_AVG = "0b100";
    parameter PRE_ITERCNT = "0b100";
    parameter PRE_RXEQ_TIMER = "0b00010100";
    parameter PRE_STEP = "STEP_SIZE_2";
    parameter PRESET_COUNT_INI = "0b0000";
    parameter PRESET_EN_LPBK_MASTER = "OTHERWISE";
    parameter PRESET_EN_LPBK_SLAVE = "OTHERWISE";
    parameter PRESET_ENABLE = "NORMAL_OP";
    parameter PRESET_EQTX_FORCE = "0b0000";
    parameter PRESET_LPBK_MASTER = "0b0000";
    parameter PRESET_LPBK_SLAVE_0 = "OTHERWISE";
    parameter PRESET_LPBK_SLAVE_1 = "OTHERWISE";
    parameter PRESET_LPBK_SLAVE_2 = "OTHERWISE";
    parameter PRESET_LPBK_SLAVE_3 = "OTHERWISE";
    parameter PRESET_REJECT = "0b00000000000";
    parameter PRESET0_POSTCURSOR = "0b1000";
    parameter PRESET0_PRECURSOR = "0b0000";
    parameter PRESET1_POSTCURSOR = "0b0101";
    parameter PRESET1_PRECURSOR = "0b0000";
    parameter PRESET10_POSTCURSOR = "0b1010";
    parameter PRESET10_PRECURSOR = "0b0000";
    parameter PRESET2_POSTCURSOR = "0b0110";
    parameter PRESET2_PRECURSOR = "0b0000";
    parameter PRESET3_POSTCURSOR = "0b0100";
    parameter PRESET3_PRECURSOR = "0b0000";
    parameter PRESET4_POSTCURSOR = "0b0000";
    parameter PRESET4_PRECURSOR = "0b0000";
    parameter PRESET5_POSTCURSOR = "0b0000";
    parameter PRESET5_PRECURSOR = "0b0011";
    parameter PRESET6_POSTCURSOR = "0b0000";
    parameter PRESET6_PRECURSOR = "0b0100";
    parameter PRESET7_POSTCURSOR = "0b0110";
    parameter PRESET7_PRECURSOR = "0b0011";
    parameter PRESET8_POSTCURSOR = "0b0100";
    parameter PRESET8_PRECURSOR = "0b0100";
    parameter PRESET9_POSTCURSOR = "0b0000";
    parameter PRESET9_PRECURSOR = "0b0101";
    parameter PS_REENTRY_TIME = "0b00000000";
    parameter RATE = "2P5G";
    parameter RATE_ENABLE = "INITIAL_SPEED_CHANGES";
    parameter RCB = "DISABLED";
    parameter REC_SPD_INFER_EQ_PH0123 = "EXCLUDE_TIME_SPENT";
    parameter REC_SPD_INFER_RCVR_CFG = "EXCLUDE_TIME_SPENT";
    parameter REC_SPD_INFER_RCVR_LOCK = "EXCLUDE_TIME_SPENT";
    parameter DIS_FUNC_B = "ENABLED";
    parameter DIS_FUNC_C = "ENABLED";
    parameter DIS_FUNC_D = "ENABLED";
    parameter REDUCE_TIMEOUTS_LTSSMSIM = "DISABLED";
    parameter REDUCE_TIMEOUTS_SIM = "DISABLED";
    parameter REDUCE_TS1 = "DISABLED";
    parameter REENTRY_DISABLE = "ENABLED";
    parameter REENTRY_TIME = "0b00000000000000";
    parameter REQ_FEEDBACK = "0b00000000";
    parameter RESET_EIEOS_INTERVAL_COUNT = "DISABLED";
    parameter REVISION_ID_ID3A = "0b00000100";
    parameter REVISION_ID_ID3B = "0b00000100";
    parameter REVISION_ID_ID3C = "0b00000100";
    parameter REVISION_ID_ID3D = "0b00000100";
    parameter RL1 = "0b0011";
    parameter RL2 = "0b0101";
    parameter RL3 = "0b0011";
    parameter ROUTING_SUPPORTED = "DISABLED";
    parameter RP_COMPLETER_EN = "DISABLED";
    parameter RSTCDR_ERR = "ENABLED";
    parameter RSTCDR_FRQ = "ENABLED";
    parameter RSTCDR_IDL = "DISABLED";
    parameter RX_BYPASS_DECODE_EN = "ENABLED";
    parameter RX_BYPASS_MSG_DEC = "NORMAL_OPERATION";
    parameter RX_CONVERT_UR_TO_CA = "NORMAL_OPERATION";
    parameter RX_D_ALLOC_C = "0b0000000001100000";
    parameter RX_D_ALLOC_N = "0b0000000000000110";
    parameter RX_D_ALLOC_P = "0b0000000001101100";
    parameter RX_DIV_MODE1 = "0b10";
    parameter RX_DIV_MODE0 = "DIV_2";
    parameter RX_DIV_MODE2 = "0b00";
    parameter RX_DL_ACTIVE_DISABLE = "BLOCK_RECEPTION_TLP";
    parameter RX_EARLY_FORWARD_DISABLE = "FWD_RX_DATA_LL";
    parameter RX_ERR_COR = "DISABLED";
    parameter RX_ERR_UCOR = "DISABLED";
    parameter RX_FORCE_RO = "DISABLED";
    parameter RX_H_ALLOC_C = "0b000000100000";
    parameter RX_H_ALLOC_N = "0b000000001000";
    parameter RX_H_ALLOC_P = "0b000000010000";
    parameter RX_HIZ = "IGNORED";
    parameter RX_IMPED_RATIO = "0b10000000";
    parameter RX_INHIBIT_ACK_NAK = "PROCESS_RCVD_ACK";
    parameter RX_INHIBIT_TLP = "PROCESS_RCVD_TLP";
    parameter RX_LCRC_INJECT_EN = "DO_NOT_INJECT_ERROR";
    parameter RX_MALF_INJECT_EN = "DO_NOT_INJECT_ERROR";
    parameter RX_POLINV = "NORMAL";
    parameter RX_PRIORITY = "DISABLED";
    parameter RX_PRIORITY_N_STARVE_THRESH = "0b00010000";
    parameter RX_PRIORITY_P_STARVE_THRESH = "0b00010000";
    parameter RX_PWRDN = "IGNORED";
    parameter RX_TLP_VALID = "DISABLED";
    parameter RXEQ_ALGO = "0b111";
    parameter RXEQ_ENABLE = "0b100";
    parameter RXEQ_EVAL_MAX = "0b11111111";
    parameter RXEQ_MANUAL = "DISABLED";
    parameter RXEQ_STATE = "0b0000";
    parameter RXF_A = "0b0100";
    parameter RXF_B = "0b0100";
    parameter RXF_C = "0b0100";
    parameter RXHF_CLKDN = "ENABLED";
    parameter RXIDLE_MAX = "0b1111";
    parameter RXIDLE_MAX2 = "0b0000010000000000";
    parameter RXIDLE_MSB = "0b11";
    parameter RXM_A = "0b10";
    parameter RXM_B = "0b01";
    parameter RXM_C = "0b00";
    parameter RXN_A = "0b00100";
    parameter RXN_B = "0b01001";
    parameter RXN_C = "0b01111";
    parameter RXOFF_SETTLE_MAX = "0b011";
    parameter RXOFF_STABLE_MAX = "0b10000";
    parameter RXPLLINIT = "DISABLED";
    parameter RXPLLRST = "SET";
    parameter SELECT_DIR_FOM_N = "FME_METHOD";
    parameter SELECTABLE_DEEMPHASIS = "6P0DB";
    parameter SEQ_NUM = "0b000000000000";
    parameter SIGNAL_DETECT_THRESHOLD = "125_MV";
    parameter SIZE_CFG0_A = "0b00000";
    parameter SIZE_CFG0_B = "0b00000";
    parameter SIZE_CFG0_C = "0b00000";
    parameter SIZE_CFG0_D = "0b00000";
    parameter SIZE_CFG1_A = "0b00000";
    parameter SIZE_CFG1_B = "0b00000";
    parameter SIZE_CFG1_C = "0b00000";
    parameter SIZE_CFG1_D = "0b00000";
    parameter SIZE_CFG2_A = "0b00000";
    parameter SIZE_CFG2_B = "0b00000";
    parameter SIZE_CFG2_C = "0b00000";
    parameter SIZE_CFG2_D = "0b00000";
    parameter SIZE_CFG3_A = "0b00000";
    parameter SIZE_CFG3_B = "0b00000";
    parameter SIZE_CFG3_C = "0b00000";
    parameter SIZE_CFG3_D = "0b00000";
    parameter SIZE_CFG4_A = "0b00000";
    parameter SIZE_CFG4_B = "0b00000";
    parameter SIZE_CFG4_C = "0b00000";
    parameter SIZE_CFG4_D = "0b00000";
    parameter SIZE_CFG5_A = "0b00000";
    parameter SIZE_CFG5_B = "0b00000";
    parameter SIZE_CFG5_C = "0b00000";
    parameter SIZE_CFG5_D = "0b00000";
    parameter SKIP_FINAL_COEF_CHECK = "DISABLED";
    parameter SLOT_CLOCK_CONFIGURATION = "REFCLK_BY_SLOT";
    parameter SLOT_IMPLEMENTED = "UNCONNECTED";
    parameter SLOT_POWER_LIMIT_SCALE = "0b00";
    parameter SLOT_POWER_LIMIT_VALUE = "0b00001010";
    parameter SPEED_LPBK_CTRL = "2P5G";
    parameter START_PRESET = "PRESET_VALUE";
    parameter START_REMOTE_ADV = "OTHERWISE";
    parameter STATE_DATA_N = "USE_RX_DATA_OBSERVATION";
    parameter STEP_SELECT = "0b00000";
    parameter STP_OVERRIDE_EN = "DISABLED";
    parameter STP_OVERRIDE_LEN = "0b00000000000";
    parameter STP_OVERRIDE_NEW_LEN = "0b00000000000";
    parameter SUBSTATE_MAX = "0b00000";
    parameter SUBSYSTEM_ID_ID2A = "0b1110000000000100";
    parameter SUBSYSTEM_ID_ID2B = "0b1110000000000100";
    parameter SUBSYSTEM_ID_ID2C = "0b1110000000000100";
    parameter SUBSYSTEM_ID_ID2D = "0b1110000000000100";
    parameter SUBSYSTEM_VENDOR_ID_ID2A = "0b0001100110101010";
    parameter SUBSYSTEM_VENDOR_ID_ID2B = "0b0001100110101010";
    parameter SUBSYSTEM_VENDOR_ID_ID2C = "0b0001100110101010";
    parameter SUBSYSTEM_VENDOR_ID_ID2D = "0b0001100110101010";
    parameter SUPP_SIZE_CFG0_A = "0b00000000000000001111";
    parameter SUPP_SIZE_CFG0_B = "0b00000000000000001111";
    parameter SUPP_SIZE_CFG0_C = "0b00000000000000001111";
    parameter SUPP_SIZE_CFG0_D = "0b00000000000000001111";
    parameter SUPP_SIZE_CFG1_A = "0b00000000000000000000";
    parameter SUPP_SIZE_CFG1_B = "0b00000000000000000000";
    parameter SUPP_SIZE_CFG1_C = "0b00000000000000000000";
    parameter SUPP_SIZE_CFG1_D = "0b00000000000000000000";
    parameter SUPP_SIZE_CFG2_A = "0b00000000000000000000";
    parameter SUPP_SIZE_CFG2_B = "0b00000000000000000000";
    parameter SUPP_SIZE_CFG2_C = "0b00000000000000000000";
    parameter SUPP_SIZE_CFG2_D = "0b00000000000000000000";
    parameter SUPP_SIZE_CFG3_A = "0b00000000000000000000";
    parameter SUPP_SIZE_CFG3_B = "0b00000000000000000000";
    parameter SUPP_SIZE_CFG3_C = "0b00000000000000000000";
    parameter SUPP_SIZE_CFG3_D = "0b00000000000000000000";
    parameter SUPP_SIZE_CFG4_A = "0b00000000000000000000";
    parameter SUPP_SIZE_CFG4_B = "0b00000000000000000000";
    parameter SUPP_SIZE_CFG4_C = "0b00000000000000000000";
    parameter SUPP_SIZE_CFG4_D = "0b00000000000000000000";
    parameter SUPP_SIZE_CFG5_A = "0b00000000000000000000";
    parameter SUPP_SIZE_CFG5_B = "0b00000000000000000000";
    parameter SUPP_SIZE_CFG5_C = "0b00000000000000000000";
    parameter SUPP_SIZE_CFG5_D = "0b00000000000000000000";
    parameter SYS_ALLOC = "PWR_BUDGET_CAP_VALUES";
    parameter T0_RX_BYPASS_MSG_DEC = "NORMAL_OPERATION";
    parameter TABLE_SIZE_MSIXCAP_A = "0b00000000111";
    parameter TABLE_SIZE_MSIXCAP_B = "0b00000000111";
    parameter TABLE_SIZE_MSIXCAP_C = "0b00000000111";
    parameter TABLE_SIZE_MSIXCAP_D = "0b00000000111";
    parameter TARGET_LINK_SPEED = "8G";
    parameter TARGET_ONLY = "DISABLED";
    parameter TD1_MEANS_ADD_HAS_N = "ECRC_CONTAINED";
    parameter TIMEOUT_THRESHOLD_PME = "0b000000000000";
    parameter TIMEOUT_THRESHOLD_PME_TO_ACK_DS = "0b00000000";
    parameter TIMER = "0b00000000";
    parameter TLP_LCRC_ERR_ENABLE = "DISABLED";
    parameter TLP_LCRC_ERR_RATE = "0b000";
    parameter TLP_SEQ_ERR_ENABLE = "DISABLED";
    parameter TLUNIT = "1_MS";
    parameter TO_EXTEND = "0b01111111";
    parameter TRNG_A0COEF = "0b101";
    parameter TRNG_A1COEF = "0b101";
    parameter TRNG_A2COEF = "0b101";
    parameter TRNG_FAST = "DISABLED";
    parameter TRNG_ITERCNT = "0b100";
    parameter TRNG_RXEQ_TIMER = "0b00100000";
    parameter TS1_ACK_BLOCK_USE_PRESET = "FORCED_TO_ZERO";
    parameter TS1_ACK_DELAY = "0b00011111";
    parameter TS1_ACK_MASK_USE_PRESET = "IGNORES_USE_PRESET";
    parameter TX_AMP_RATIO_MARGIN0_FULL = "0b10000000";
    parameter TX_AMP_RATIO_MARGIN0_HALF = "0b01010000";
    parameter TX_AMP_RATIO_MARGIN1_FULL = "0b01111000";
    parameter TX_AMP_RATIO_MARGIN1_HALF = "0b01011000";
    parameter TX_AMP_RATIO_MARGIN2_FULL = "0b01101000";
    parameter TX_AMP_RATIO_MARGIN2_HALF = "0b01001000";
    parameter TX_AMP_RATIO_MARGIN3_FULL = "0b01100000";
    parameter TX_AMP_RATIO_MARGIN3_HALF = "0b01000000";
    parameter TX_AMP_RATIO_MARGIN4_FULL = "0b01011000";
    parameter TX_AMP_RATIO_MARGIN4_HALF = "0b00111000";
    parameter TX_AMP_RATIO_MARGIN5_FULL = "0b01010000";
    parameter TX_AMP_RATIO_MARGIN5_HALF = "0b00110000";
    parameter TX_AMP_RATIO_MARGIN6_FULL = "0b01001000";
    parameter TX_AMP_RATIO_MARGIN6_HALF = "0b00101000";
    parameter TX_AMP_RATIO_MARGIN7_FULL = "0b01000000";
    parameter TX_AMP_RATIO_MARGIN7_HALF = "0b00100000";
    parameter TX_BYPASS_DECODE_EN = "ENABLED";
    parameter TX_BYPASS_MSG_DEC = "NORMAL_OPERATION";
    parameter TX_COMP_RECEIVE = "DOES_NOT_ASSERT";
    parameter TX_CONVERT_UR_TO_CA = "NORMAL_OPERATION";
    parameter TX_D_ALLOC_C = "0b0000000001100000";
    parameter TX_D_ALLOC_N = "0b0000000000000110";
    parameter TX_D_ALLOC_P = "0b0000000001101100";
    parameter TX_DIV_MODE0 = "0b10";
    parameter TX_DIV_MODE1 = "0b10";
    parameter TX_DIV_MODE2 = "0b10";
    parameter TX_EQ_EVAL_CNT_SEL = "WAIT_8_CLKS";
    parameter TX_ERR_COR = "DISABLED";
    parameter TX_ERR_UCOR = "DISABLED";
    parameter TX_FORCE_RO = "DISABLED";
    parameter TX_GAP_INJECT_EN = "DO_NOT_INJECT_GAP";
    parameter TX_H_ALLOC_C = "0b000000100000";
    parameter TX_H_ALLOC_N = "0b000000001000";
    parameter TX_H_ALLOC_P = "0b000000010000";
    parameter TX_HIZ = "IGNORED";
    parameter TX_IMPED_RATIO = "0b10000000";
    parameter TX_PAR1_INJECT_EN = "DO_NOT_INJECT_ERR";
    parameter TX_PAR2_HANDLE_DISABLE = "ENABLE_HANDLING";
    parameter TX_PAR2_INJECT_EN = "DO_NOT_INJECT_ERR";
    parameter TX_PAR2_REPORT_DISABLE = "ENABLE_REPORTING";
    parameter TX_POLINV = "NORMAL";
    parameter TX_PRE_RATIO = "0b00000000";
    parameter TX_PRE_RATIO_DEEMP0_FULL = "0b00000000";
    parameter TX_PRE_RATIO_DEEMP0_HALF = "0b00000000";
    parameter TX_PRE_RATIO_DEEMP1_FULL = "0b00000000";
    parameter TX_PRE_RATIO_DEEMP1_HALF = "0b00000000";
    parameter TX_PRIORITY = "DISABLED";
    parameter TX_PRIORITY_N_STARVE_THRESH = "0b00010000";
    parameter TX_PRIORITY_P_STARVE_THRESH = "0b00010000";
    parameter TX_PST_RATIO = "0b00010101";
    parameter TX_PST_RATIO_DEEMP0_FULL = "0b00100000";
    parameter TX_PST_RATIO_DEEMP0_HALF = "0b00100000";
    parameter TX_PST_RATIO_DEEMP1_FULL = "0b00010101";
    parameter TX_PST_RATIO_DEEMP1_HALF = "0b00010101";
    parameter TX_QUIESCE = "DISABLED";
    parameter TX_REPLAY_ECC1_HANDLE_DISABLE = "ENABLE_CORRECTION";
    parameter TX_REPLAY_ECC1_INJECT_EN = "DO_NOT_INJECT_ERR";
    parameter TX_REPLAY_ECC1_REPORT_DISABLE = "ENABLE_REPORTING";
    parameter TX_REPLAY_ECC2_HANDLE_DISABLE = "ENABLE_HANDLING";
    parameter TX_REPLAY_ECC2_INJECT_EN = "DO_NOT_INJECT_ERR";
    parameter TX_REPLAY_ECC2_REPORT_DISABLE = "ENABLE_REPORTING";
    parameter TX_REQ_EQ = "DISABLED";
    parameter TX_SELECT_RX_FEEDBACK = "REFCLK";
    parameter TX_TLP_VALID = "DISABLED";
    parameter TXF_A = "0b0100";
    parameter TXF_B = "0b0100";
    parameter TXF_C = "0b0100";
    parameter TXHF_CLKDN = "ENABLED";
    parameter TXM_A = "0b10";
    parameter TXM_B = "0b01";
    parameter TXM_C = "0b00";
    parameter TXN_A = "0b00100";
    parameter TXN_B = "0b01001";
    parameter TXN_C = "0b01111";
    parameter TXPLL_INIT = "DISABLED";
    parameter TXPLLRST = "DISABLED";
    parameter TYPE1_TYPE0_N = "ENDPOINT";
    parameter U_CLK_PERIOD = "0b0001111101000000";
    parameter US_PORT_PS_ENTRY_TIME = "0b0000000000000000";
    parameter US_PORT_RX_PRESET_HINT = "0b010";
    parameter US_PORT_TX_PRESET = "0b0100";
    parameter USE_COEF_PRE_MTHD_CTRL = "PRESET_VALUE";
    parameter USE_COEF_UPDN_CTRL = "PRESET_VALUE";
    parameter USER_AUTO_N = "AUTOMATIC_ON_RECEPTION";
    parameter VEC_MASK_CAPABLE_MSICAP_A = "ENABLED";
    parameter VEC_MASK_CAPABLE_MSICAP_B = "ENABLED";
    parameter VEC_MASK_CAPABLE_MSICAP_C = "ENABLED";
    parameter VEC_MASK_CAPABLE_MSICAP_D = "ENABLED";
    parameter VENDOR_ID_ID1A = "0b0001100110101010";
    parameter VENDOR_ID_ID1B = "0b0001100110101010";
    parameter VENDOR_ID_ID1C = "0b0001100110101010";
    parameter VENDOR_ID_ID1D = "0b0001100110101010";
    parameter VENDOR0_UR = "REPORT";
    parameter VERSION_AER_CAP = "VER_0X2";
    parameter VERSION_PM_CAP = "0b011";
    parameter XLCY0 = "0b00000000";
    parameter XLCY1 = "0b00000000";
    parameter RX_ESP_RESP_WAIT = "0b01000000";
    parameter SEL_PCLK_DIV2 = "PCLK_DIV2";
    parameter COMPLIANCE = "ENABLED";
    parameter LOOPBACK = "ENABLED";
    parameter HOT_RESET = "ENABLED";
    parameter DIS_PREVENT = "ENABLED";
    parameter MPS_VIOLATION_RX = "DISABLED";
    parameter MPS_VIOLATION_TX = "DISABLED";
    parameter EN_RX_ALLOC_SEL = "HW";
    parameter EN_TX_ALLOC_SEL = "HW";
    parameter AUX_CLK_PERIOD = "0b1111010000100100";
    parameter EN_PIPE_IF_CTRL = "DISABLED";
    parameter PIPE_PWRDN = "P1";
    parameter TX_CM_DIS = "DEASSERTED";
    parameter RX_EI_DIS = "DEASSERTED";
    parameter PCLKREQ_N = "DEASSERTED";
    parameter STS_PHY_STATUS = "DEASSERTED";
    parameter STS_PIPE_RSTN = "DEASSERTED";
    parameter LEGACY_MODE = "MATCH_TS";
    parameter OVERFLOW = "DISABLED";
    parameter DIR = "RECEIVE";
    parameter SPEED = "8G";
    parameter LANE = "0";
    parameter COEF_ENABLE_8G = "DISABLED";
    parameter PRESET_ENABLE_8G = "DISABLED";
    parameter VALUE_8G_PRE = "0b000000";
    parameter VALUE_8G_POST = "0b000000";
    parameter REQ_EQ_MAX_COUNT = "0b10";
    parameter MESO_LPBK = "DISABLED";
    parameter TX_REPLAY_ECC2_INJECT_M_1_N = "INJECT_1_ERR";
    parameter TX_REPLAY_ECC1_INJECT_M_1_N = "INJECT_1_ERR";
    parameter REDO = "DISABLED";
    parameter RX_PAR_REPORT_DISABLE = "ENABLE_REPORTING";
    parameter RX_PAR_INJECT_EN = "DO_NOT_INJECT_ERR";
    parameter RX_ECC2_REPORT_DISABLE = "ENABLE_REPORTING";
    parameter RX_ECC2_HANDLE_DISABLE = "ENABLE_HANDLING";
    parameter RX_ECC2_INJECT_M_1_N = "INJECT_1_ERR";
    parameter RX_ECC2_INJECT_TYPE = "POSTED_DATA_RAM";
    parameter RX_ECC2_INJECT_EN = "DO_NOT_INJECT_ERR";
    parameter RX_ECC1_REPORT_DISABLE = "ENABLE_REPORTING";
    parameter RX_ECC1_HANDLE_DISABLE = "ENABLE_HANDLING";
    parameter RX_ECC1_INJECT_M_1_N = "INJECT_1_ERR";
    parameter RX_ECC1_INJECT_TYPE = "POSTED_DATA_RAM";
    parameter RX_ECC1_INJECT_EN = "DO_NOT_INJECT_ERR";
    parameter RX_ERR_PAR = "OTHERWISE";
    parameter RX_ERR_ECC2 = "OTHERWISE";
    parameter RX_ERR_ECC1 = "OTHERWISE";
    parameter TX_PAR_REPORT_DISABLE = "ENABLE_REPORTING";
    parameter TX_PAR_INJECT_EN = "DO_NOT_INJECT_ERR";
    parameter TX_ECC2_REPORT_DISABLE = "ENABLE_REPORTING";
    parameter TX_ECC2_HANDLE_DISABLE = "ENABLE_HANDLING";
    parameter TX_ECC2_INJECT_M_1_N = "INJECT_1_ERR";
    parameter TX_ECC2_INJECT_TYPE = "POSTED_DATA_RAM";
    parameter TX_ECC2_INJECT_EN = "DO_NOT_INJECT_ERR";
    parameter TX_ECC1_REPORT_DISABLE = "ENABLE_REPORTING";
    parameter TX_ECC1_HANDLE_DISABLE = "ENABLE_HANDLING";
    parameter TX_ECC1_INJECT_M_1_N = "INJECT_1_ERR";
    parameter TX_ECC1_INJECT_TYPE = "POSTED_DATA_RAM";
    parameter TX_ECC1_INJECT_EN = "DO_NOT_INJECT_ERR";
    parameter TX_ERR_PAR = "OTHERWISE";
    parameter TX_ERR_ECC2 = "OTHERWISE";
    parameter TX_ERR_ECC1 = "OTHERWISE";
    parameter MAX_PAYLOAD_SIZE_SUPPORTED = "256_BYTES";
    parameter ARXCAL_OUT = "DISABLED";
    parameter F_ARXDPDIR = "IGNORED";
    parameter IDLE_INFER_REC_RCVR_CFG = "OTHERWISE";
    parameter IDLE_INFER_LPBK_SLAVE = "OTHERWISE";
    parameter IDLE_INFER_REC_SPEED2_SUCCESS = "OTHERWISE";
    parameter IDLE_INFER_REC_SPEED2_UNSUCCESS = "OTHERWISE";
    parameter IDLE_INFER_L0_TO_REC_RCVR_LOCK = "OTHERWISE";
    parameter SPEED_CHANGE_FAIL = "OTHERWISE";
    parameter DIRECT_TO_DETECT_FAST = "OTHERWISE";
    parameter DIRECT_TO_RCVRY_CH_BOND = "OTHERWISE";
    parameter DIRECT_TO_LPBK_ENTRY = "OTHERWISE";
    parameter DIRECT_SPEED_CHANGE = "OTHERWISE";
    parameter L0_TO_REC_RCVR_LOCK_RX_TS12 = "OTHERWISE";
    parameter L0_TO_REC_RCVR_LOCK_RX_8G_EIE = "OTHERWISE";
    parameter L0_TO_REC_RCVR_LOCK_RX_INFER = "OTHERWISE";
    parameter DIRECT_TO_RCVRY_PHY = "OTHERWISE";
    parameter DIRECT_TO_RCVRY_FRAME = "OTHERWISE";
    parameter DIRECT_TO_RCVRY_REPLAY = "OTHERWISE";
    parameter DIRECT_TO_HOT_RESET = "OTHERWISE";
    parameter DIRECT_TO_DISABLE = "OTHERWISE";
    parameter RX_L0S_DIRECT_TO_RCVRY = "OTHERWISE";
    parameter AUTONOMOUS_WIDTH_CHANGE = "OTHERWISE";
    parameter DIRECTED_RETRAIN_LINK = "OTHERWISE";
    parameter ERR_TX_PIPE_UNDERFLOW = "OTHERWISE";
    parameter TS2_DETECT3 = "OTHERWISE";
    parameter TS2_DETECT2 = "OTHERWISE";
    parameter TS2_DETECT1 = "OTHERWISE";
    parameter TS2_DETECT0 = "OTHERWISE";
    parameter TS1_DETECT3 = "OTHERWISE";
    parameter TS1_DETECT2 = "OTHERWISE";
    parameter TS1_DETECT1 = "OTHERWISE";
    parameter TS1_DETECT0 = "OTHERWISE";
    parameter TS2I_DETECT3 = "OTHERWISE";
    parameter TS2I_DETECT2 = "OTHERWISE";
    parameter TS2I_DETECT1 = "OTHERWISE";
    parameter TS2I_DETECT0 = "OTHERWISE";
    parameter TS1I_DETECT3 = "OTHERWISE";
    parameter TS1I_DETECT2 = "OTHERWISE";
    parameter TS1I_DETECT1 = "OTHERWISE";
    parameter TS1I_DETECT0 = "OTHERWISE";
    parameter FTS_DETECT3 = "OTHERWISE";
    parameter FTS_DETECT2 = "OTHERWISE";
    parameter FTS_DETECT1 = "OTHERWISE";
    parameter FTS_DETECT0 = "OTHERWISE";
    parameter SKP_DETECT3 = "OTHERWISE";
    parameter SKP_DETECT2 = "OTHERWISE";
    parameter SKP_DETECT1 = "OTHERWISE";
    parameter SKP_DETECT0 = "OTHERWISE";
    parameter EIE_DETECT3 = "OTHERWISE";
    parameter EIE_DETECT2 = "OTHERWISE";
    parameter EIE_DETECT1 = "OTHERWISE";
    parameter EIE_DETECT0 = "OTHERWISE";
    parameter EIOS_DETECT3 = "OTHERWISE";
    parameter EIOS_DETECT2 = "OTHERWISE";
    parameter EIOS_DETECT1 = "OTHERWISE";
    parameter EIOS_DETECT0 = "OTHERWISE";
    parameter DATA_DETECT3 = "OTHERWISE";
    parameter DATA_DETECT2 = "OTHERWISE";
    parameter DATA_DETECT1 = "OTHERWISE";
    parameter DATA_DETECT0 = "OTHERWISE";
    parameter SDS_DETECT3 = "OTHERWISE";
    parameter SDS_DETECT2 = "OTHERWISE";
    parameter SDS_DETECT1 = "OTHERWISE";
    parameter SDS_DETECT0 = "OTHERWISE";
    parameter INFO_BAD_TLP_NULL_ERR = "OTHERWISE";
    parameter INFO_BAD_TLP_PHY_ERR = "OTHERWISE";
    parameter INFO_BAD_TLP_MALF_ERR = "OTHERWISE";
    parameter INFO_BAD_TLP_ECRC_ERR = "OTHERWISE";
    parameter INFO_SCHEDULE_DUPL_ACK = "OTHERWISE";
    parameter INFO_BAD_TLP_SEQ_ERR = "OTHERWISE";
    parameter INFO_BAD_TLP_CRC_ERR = "OTHERWISE";
    parameter INFO_NAK_RECEIVED = "OTHERWISE";
    parameter INFO_DESKEW_OVERFLOW_ERROR = "OTHERWISE";
    parameter INFO_TX_DATA_UNDERFLOW = "OTHERWISE";
    parameter INFO_REPLAY_STARTED = "OTHERWISE";
    parameter ERR_AER_TX_PAR2 = "OTHERWISE";
    parameter ERR_AER_TX_REPLAY_ECC2 = "OTHERWISE";
    parameter ERR_AER_TX_REPLAY_ECC1 = "OTHERWISE";
    parameter ERR_AER_SURPRISE_DOWN = "OTHERWISE";
    parameter ERR_AER_DL_PROTOCOL_ERROR = "OTHERWISE";
    parameter ERR_AER_REPLAY_TIMER_TIMEOUT = "OTHERWISE";
    parameter ERR_AER_REPLAY_NUM_ROLLOVER = "OTHERWISE";
    parameter ERR_AER_BAD_DLLP = "OTHERWISE";
    parameter ERR_AER_BAD_TLP = "OTHERWISE";
    parameter ERR_AER_RECEIVER_ERROR = "OTHERWISE";
    parameter P_RX_LIM_H = "DISABLED";
    parameter P_RX_LIM_D = "DISABLED";
    parameter N_RX_LIM_H = "DISABLED";
    parameter N_RX_LIM_D = "DISABLED";
    parameter C_RX_LIM_H = "DISABLED";
    parameter C_RX_LIM_D = "DISABLED";
    parameter P_TX_LIM_H = "DISABLED";
    parameter P_TX_LIM_D = "DISABLED";
    parameter N_TX_LIM_H = "DISABLED";
    parameter N_TX_LIM_D = "DISABLED";
    parameter C_TX_LIM_H = "DISABLED";
    parameter C_TX_LIM_D = "DISABLED";
    parameter MAX_RSA_WAIT = "0b00101000";
    parameter F_ARXDPNULL = "0b00000";
endmodule

module PDP16K_MODE(DI0, DI1, DI2, DI3, DI4, DI5, DI6, DI7, DI8, DI9, DI10, DI11, DI12, DI13, DI14, DI15, DI16, DI17, DI18, DI19, DI20, DI21, DI22, DI23, DI24, DI25, DI26, DI27, DI28, DI29, DI30, DI31, DI32, DI33, DI34, DI35, ADW0, ADW1, ADW2, ADW3, ADW4, ADW5, ADW6, ADW7, ADW8, ADW9, ADW10, ADW11, ADW12, ADW13, ADR0, ADR1, ADR2, ADR3, ADR4, ADR5, ADR6, ADR7, ADR8, ADR9, ADR10, ADR11, ADR12, ADR13, CLKW, CLKR, CEW, CER, CSW0, CSW1, CSW2, CSR0, CSR1, CSR2, RST, DO0, DO1, DO2, DO3, DO4, DO5, DO6, DO7, DO8, DO9, DO10, DO11, DO12, DO13, DO14, DO15, DO16, DO17, DO18, DO19, DO20, DO21, DO22, DO23, DO24, DO25, DO26, DO27, DO28, DO29, DO30, DO31, DO32, DO33, DO34, DO35, ONEBITERR, TWOBITERR); //synthesis syn_black_box syn_lib_cell=1
    input DI0;
    input DI1;
    input DI2;
    input DI3;
    input DI4;
    input DI5;
    input DI6;
    input DI7;
    input DI8;
    input DI9;
    input DI10;
    input DI11;
    input DI12;
    input DI13;
    input DI14;
    input DI15;
    input DI16;
    input DI17;
    input DI18;
    input DI19;
    input DI20;
    input DI21;
    input DI22;
    input DI23;
    input DI24;
    input DI25;
    input DI26;
    input DI27;
    input DI28;
    input DI29;
    input DI30;
    input DI31;
    input DI32;
    input DI33;
    input DI34;
    input DI35;
    input ADW0;
    input ADW1;
    input ADW2;
    input ADW3;
    input ADW4;
    input ADW5;
    input ADW6;
    input ADW7;
    input ADW8;
    input ADW9;
    input ADW10;
    input ADW11;
    input ADW12;
    input ADW13;
    input ADR0;
    input ADR1;
    input ADR2;
    input ADR3;
    input ADR4;
    input ADR5;
    input ADR6;
    input ADR7;
    input ADR8;
    input ADR9;
    input ADR10;
    input ADR11;
    input ADR12;
    input ADR13;
    input CLKW;
    input CLKR;
    input CEW;
    input CER;
    input CSW0;
    input CSW1;
    input CSW2;
    input CSR0;
    input CSR1;
    input CSR2;
    input RST;
    output DO0;
    output DO1;
    output DO2;
    output DO3;
    output DO4;
    output DO5;
    output DO6;
    output DO7;
    output DO8;
    output DO9;
    output DO10;
    output DO11;
    output DO12;
    output DO13;
    output DO14;
    output DO15;
    output DO16;
    output DO17;
    output DO18;
    output DO19;
    output DO20;
    output DO21;
    output DO22;
    output DO23;
    output DO24;
    output DO25;
    output DO26;
    output DO27;
    output DO28;
    output DO29;
    output DO30;
    output DO31;
    output DO32;
    output DO33;
    output DO34;
    output DO35;
    output ONEBITERR;
    output TWOBITERR;
    parameter DATA_WIDTH_W = "X36";
    parameter DATA_WIDTH_R = "X36";
    parameter OUTREG = "BYPASSED";
    parameter RESETMODE = "SYNC";
    parameter GSR = "ENABLED";
    parameter ECC = "DISABLED";
    parameter INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter CSDECODE_W = "000";
    parameter CSDECODE_R = "000";
    parameter ASYNC_RST_RELEASE = "SYNC";
    parameter INIT_DATA = "STATIC";
endmodule

module PDP16K(DI, ADW, ADR, CLKW, CLKR, CEW, CER, CSW, CSR, RST, DO, ONEBITERR, TWOBITERR); //synthesis syn_black_box syn_lib_cell=1
    input [35:0] DI;
    input [13:0] ADW;
    input [13:0] ADR;
    input CLKW;
    input CLKR;
    input CEW;
    input CER;
    input [2:0] CSW;
    input [2:0] CSR;
    input RST;
    output [35:0] DO;
    output ONEBITERR;
    output TWOBITERR;
    parameter DATA_WIDTH_W = "X36";
    parameter DATA_WIDTH_R = "X36";
    parameter OUTREG = "BYPASSED";
    parameter RESETMODE = "SYNC";
    parameter GSR = "ENABLED";
    parameter ECC = "DISABLED";
    parameter INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter CSDECODE_W = "000";
    parameter CSDECODE_R = "000";
    parameter ASYNC_RST_RELEASE = "SYNC";
    parameter INIT_DATA = "STATIC";
endmodule

module PDPSC16K_MODE(DI0, DI1, DI2, DI3, DI4, DI5, DI6, DI7, DI8, DI9, DI10, DI11, DI12, DI13, DI14, DI15, DI16, DI17, DI18, DI19, DI20, DI21, DI22, DI23, DI24, DI25, DI26, DI27, DI28, DI29, DI30, DI31, DI32, DI33, DI34, DI35, ADW0, ADW1, ADW2, ADW3, ADW4, ADW5, ADW6, ADW7, ADW8, ADW9, ADW10, ADW11, ADW12, ADW13, ADR0, ADR1, ADR2, ADR3, ADR4, ADR5, ADR6, ADR7, ADR8, ADR9, ADR10, ADR11, ADR12, ADR13, CLK, CER, CEW, CSW0, CSW1, CSW2, CSR0, CSR1, CSR2, RST, DO0, DO1, DO2, DO3, DO4, DO5, DO6, DO7, DO8, DO9, DO10, DO11, DO12, DO13, DO14, DO15, DO16, DO17, DO18, DO19, DO20, DO21, DO22, DO23, DO24, DO25, DO26, DO27, DO28, DO29, DO30, DO31, DO32, DO33, DO34, DO35, ONEBITERR, TWOBITERR); //synthesis syn_black_box syn_lib_cell=1
    input DI0;
    input DI1;
    input DI2;
    input DI3;
    input DI4;
    input DI5;
    input DI6;
    input DI7;
    input DI8;
    input DI9;
    input DI10;
    input DI11;
    input DI12;
    input DI13;
    input DI14;
    input DI15;
    input DI16;
    input DI17;
    input DI18;
    input DI19;
    input DI20;
    input DI21;
    input DI22;
    input DI23;
    input DI24;
    input DI25;
    input DI26;
    input DI27;
    input DI28;
    input DI29;
    input DI30;
    input DI31;
    input DI32;
    input DI33;
    input DI34;
    input DI35;
    input ADW0;
    input ADW1;
    input ADW2;
    input ADW3;
    input ADW4;
    input ADW5;
    input ADW6;
    input ADW7;
    input ADW8;
    input ADW9;
    input ADW10;
    input ADW11;
    input ADW12;
    input ADW13;
    input ADR0;
    input ADR1;
    input ADR2;
    input ADR3;
    input ADR4;
    input ADR5;
    input ADR6;
    input ADR7;
    input ADR8;
    input ADR9;
    input ADR10;
    input ADR11;
    input ADR12;
    input ADR13;
    input CLK;
    input CER;
    input CEW;
    input CSW0;
    input CSW1;
    input CSW2;
    input CSR0;
    input CSR1;
    input CSR2;
    input RST;
    output DO0;
    output DO1;
    output DO2;
    output DO3;
    output DO4;
    output DO5;
    output DO6;
    output DO7;
    output DO8;
    output DO9;
    output DO10;
    output DO11;
    output DO12;
    output DO13;
    output DO14;
    output DO15;
    output DO16;
    output DO17;
    output DO18;
    output DO19;
    output DO20;
    output DO21;
    output DO22;
    output DO23;
    output DO24;
    output DO25;
    output DO26;
    output DO27;
    output DO28;
    output DO29;
    output DO30;
    output DO31;
    output DO32;
    output DO33;
    output DO34;
    output DO35;
    output ONEBITERR;
    output TWOBITERR;
    parameter DATA_WIDTH_W = "X36";
    parameter DATA_WIDTH_R = "X36";
    parameter OUTREG = "BYPASSED";
    parameter RESETMODE = "SYNC";
    parameter GSR = "ENABLED";
    parameter ECC = "DISABLED";
    parameter INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter CSDECODE_W = "000";
    parameter CSDECODE_R = "000";
    parameter ASYNC_RST_RELEASE = "SYNC";
    parameter INIT_DATA = "STATIC";
endmodule

module PDPSC16K(DI, ADW, ADR, CLK, CER, CEW, CSW, CSR, RST, DO, ONEBITERR, TWOBITERR); //synthesis syn_black_box syn_lib_cell=1
    input [35:0] DI;
    input [13:0] ADW;
    input [13:0] ADR;
    input CLK;
    input CER;
    input CEW;
    input [2:0] CSW;
    input [2:0] CSR;
    input RST;
    output [35:0] DO;
    output ONEBITERR;
    output TWOBITERR;
    parameter DATA_WIDTH_W = "X36";
    parameter DATA_WIDTH_R = "X36";
    parameter OUTREG = "BYPASSED";
    parameter RESETMODE = "SYNC";
    parameter GSR = "ENABLED";
    parameter ECC = "DISABLED";
    parameter INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter CSDECODE_W = "000";
    parameter CSDECODE_R = "000";
    parameter ASYNC_RST_RELEASE = "SYNC";
    parameter INIT_DATA = "STATIC";
endmodule

module PDPSC512K(DI, ADW, ADR, CLK, CEW, CER, WE, CSW, CSR, RSTR, BYTEEN_N, DO, ERRDECA, ERRDECB); //synthesis syn_black_box syn_lib_cell=1
    input [31:0] DI;
    input [13:0] ADW;
    input [13:0] ADR;
    input CLK;
    input CEW;
    input CER;
    input WE;
    input CSW;
    input CSR;
    input RSTR;
    input [3:0] BYTEEN_N;
    output [31:0] DO;
    output [1:0] ERRDECA;
    output [1:0] ERRDECB;
    parameter OUTREG = "NO_REG";
    parameter GSR = "ENABLED";
    parameter RESETMODE = "SYNC";
    parameter INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_40 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_41 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_42 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_43 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_44 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_45 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_46 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_47 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_48 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_49 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_4A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_4B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_4C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_4D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_4E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_4F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_50 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_51 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_52 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_53 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_54 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_55 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_56 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_57 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_58 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_59 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_5A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_5B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_5C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_5D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_5E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_5F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_60 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_61 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_62 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_63 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_64 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_65 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_66 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_67 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_68 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_69 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_6A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_6B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_6C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_6D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_6E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_6F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_70 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_71 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_72 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_73 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_74 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_75 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_76 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_77 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_78 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_79 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_7A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_7B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_7C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_7D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_7E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_7F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter ASYNC_RESET_RELEASE = "SYNC";
    parameter ECC_BYTE_SEL = "ECC_EN";
endmodule


module PLL(INTFBKOP, INTFBKOS, INTFBKOS2, INTFBKOS3, INTFBKOS4, INTFBKOS5, DIR, DIRSEL, LOADREG, DYNROTATE, LMMICLK, LMMIRESET_N, LMMIREQUEST, LMMIWRRD_N, LMMIOFFSET, LMMIWDATA, LMMIRDATA, LMMIRDATAVALID, LMMIREADY, PLLPOWERDOWN_N, REFCK, CLKOP, CLKOS, CLKOS2, CLKOS3, CLKOS4, CLKOS5, ENCLKOP, ENCLKOS, ENCLKOS2, ENCLKOS3, ENCLKOS4, ENCLKOS5, FBKCK, INTLOCK, LEGACY, LEGRDYN, LOCK, PFDDN, PFDUP, PLLRESET, STDBY, REFMUXCK, REGQA, REGQB, REGQB1, CLKOUTDL, ROTDEL, DIRDEL, ROTDELP1, GRAYTEST, BINTEST, DIRDELP1, GRAYACT, BINACT); //synthesis syn_black_box syn_lib_cell=1
    output INTFBKOP;
    output INTFBKOS;
    output INTFBKOS2;
    output INTFBKOS3;
    output INTFBKOS4;
    output INTFBKOS5;
    input DIR;
    input [2:0] DIRSEL;
    input LOADREG;
    input DYNROTATE;
    input LMMICLK;
    input LMMIRESET_N;
    input LMMIREQUEST;
    input LMMIWRRD_N;
    input [6:0] LMMIOFFSET;
    input [7:0] LMMIWDATA;
    output [7:0] LMMIRDATA;
    output LMMIRDATAVALID;
    output LMMIREADY;
    input PLLPOWERDOWN_N;
    input REFCK;
    output CLKOP;
    output CLKOS;
    output CLKOS2;
    output CLKOS3;
    output CLKOS4;
    output CLKOS5;
    input ENCLKOP;
    input ENCLKOS;
    input ENCLKOS2;
    input ENCLKOS3;
    input ENCLKOS4;
    input ENCLKOS5;
    input FBKCK;
    output INTLOCK;
    input LEGACY;
    output LEGRDYN;
    output LOCK;
    output PFDDN;
    output PFDUP;
    input PLLRESET;
    input STDBY;
    output REFMUXCK;
    output REGQA;
    output REGQB;
    output REGQB1;
    output CLKOUTDL;
    input ROTDEL;
    input DIRDEL;
    input ROTDELP1;
    input [4:0] GRAYTEST;
    input [1:0] BINTEST;
    input DIRDELP1;
    input [4:0] GRAYACT;
    input [1:0] BINACT;
    parameter BW_CTL_BIAS = "0b0101";
    parameter CLKOP_TRIM = "0b0000";
    parameter CLKOS_TRIM = "0b0000";
    parameter CLKOS2_TRIM = "0b0000";
    parameter CLKOS3_TRIM = "0b0000";
    parameter CLKOS4_TRIM = "0b0000";
    parameter CLKOS5_TRIM = "0b0000";
    parameter CRIPPLE = "5P";
    parameter CSET = "40P";
    parameter DELAY_CTRL = "200PS";
    parameter DELA = "0";
    parameter DELB = "0";
    parameter DELC = "0";
    parameter DELD = "0";
    parameter DELE = "0";
    parameter DELF = "0";
    parameter DIRECTION = "DISABLED";
    parameter DIVA = "0";
    parameter DIVB = "0";
    parameter DIVC = "0";
    parameter DIVD = "0";
    parameter DIVE = "0";
    parameter DIVF = "0";
    parameter DYN_SEL = "0b000";
    parameter DYN_SOURCE = "STATIC";
    parameter ENCLK_CLKOP = "DISABLED";
    parameter ENCLK_CLKOS = "DISABLED";
    parameter ENCLK_CLKOS2 = "DISABLED";
    parameter ENCLK_CLKOS3 = "DISABLED";
    parameter ENCLK_CLKOS4 = "DISABLED";
    parameter ENCLK_CLKOS5 = "DISABLED";
    parameter ENABLE_SYNC = "DISABLED";
    parameter FAST_LOCK_EN = "ENABLED";
    parameter V2I_1V_EN = "DISABLED";
    parameter FBK_CUR_BLE = "0b00000000";
    parameter FBK_EDGE_SEL = "POSITIVE";
    parameter FBK_IF_TIMING_CTL = "0b00";
    parameter FBK_INTEGER_MODE = "DISABLED";
    parameter FBK_MASK = "0b00001000";
    parameter FBK_MMD_DIG = "8";
    parameter FBK_MMD_PULS_CTL = "0b0000";
    parameter FBK_MODE = "0b00";
    parameter FBK_PI_BYPASS = "NOT_BYPASSED";
    parameter FBK_PI_RC = "0b1100";
    parameter FBK_PR_CC = "0b0000";
    parameter FBK_PR_IC = "0b1000";
    parameter FLOAT_CP = "DISABLED";
    parameter FLOCK_CTRL = "2X";
    parameter FLOCK_EN = "ENABLED";
    parameter FLOCK_SRC_SEL = "REFCLK";
    parameter FORCE_FILTER = "DISABLED";
    parameter I_CTRL = "10UA";
    parameter IPI_CMP = "0b1000";
    parameter IPI_CMPN = "0b0011";
    parameter IPI_COMP_EN = "DISABLED";
    parameter IPP_CTRL = "0b1000";
    parameter IPP_SEL = "0b1111";
    parameter KP_VCO = "0b11001";
    parameter LDT_INT_LOCK_STICKY = "DISABLED";
    parameter LDT_LOCK = "1536CYC";
    parameter LDT_LOCK_SEL = "U_FREQ";
    parameter LEGACY_ATT = "DISABLED";
    parameter LOAD_REG = "DISABLED";
    parameter OPENLOOP_EN = "DISABLED";
    parameter PHIA = "0";
    parameter PHIB = "0";
    parameter PHIC = "0";
    parameter PHID = "0";
    parameter PHIE = "0";
    parameter PHIF = "0";
    parameter PLLPDN_EN = "DISABLED";
    parameter PLLPD_N = "UNUSED";
    parameter PLLRESET_ENA = "DISABLED";
    parameter REF_INTEGER_MODE = "DISABLED";
    parameter REF_MASK = "0b00000000";
    parameter REF_MMD_DIG = "8";
    parameter REF_MMD_IN = "0b00001000";
    parameter REF_MMD_PULS_CTL = "0b0000";
    parameter REF_TIMING_CTL = "0b00";
    parameter REFIN_RESET = "SET";
    parameter RESET_LF = "DISABLED";
    parameter ROTATE = "DISABLED";
    parameter SEL_OUTA = "DISABLED";
    parameter SEL_OUTB = "DISABLED";
    parameter SEL_OUTC = "DISABLED";
    parameter SEL_OUTD = "DISABLED";
    parameter SEL_OUTE = "DISABLED";
    parameter SEL_OUTF = "DISABLED";
    parameter SLEEP = "DISABLED";
    parameter SSC_DITHER = "DISABLED";
    parameter SSC_EN_CENTER_IN = "DOWN_TRIANGLE";
    parameter SSC_EN_SDM = "DISABLED";
    parameter SSC_EN_SSC = "DISABLED";
    parameter SSC_F_CODE = "0b000000000000000";
    parameter SSC_N_CODE = "0b000010100";
    parameter SSC_ORDER = "SDM_ORDER2";
    parameter SSC_PI_BYPASS = "NOT_BYPASSED";
    parameter SSC_REG_WEIGHTING_SEL = "0b000";
    parameter SSC_SQUARE_MODE = "DISABLED";
    parameter SSC_STEP_IN = "0b0000000";
    parameter SSC_TBASE = "0b000000000000";
    parameter STDBY_ATT = "DISABLED";
    parameter TRIMOP_BYPASS_N = "BYPASSED";
    parameter TRIMOS_BYPASS_N = "BYPASSED";
    parameter TRIMOS2_BYPASS_N = "BYPASSED";
    parameter TRIMOS3_BYPASS_N = "BYPASSED";
    parameter TRIMOS4_BYPASS_N = "BYPASSED";
    parameter TRIMOS5_BYPASS_N = "BYPASSED";
    parameter V2I_KVCO_SEL = "85";
    parameter V2I_PP_ICTRL = "0b00110";
    parameter V2I_PP_RES = "10K";
    parameter CLKMUX_FB = "CMUX_CLKOP";
    parameter SEL_FBK = "DIVA";
    parameter DIV_DEL = "0b0000001";
    parameter PHASE_SEL_DEL = "0b000";
    parameter PHASE_SEL_DEL_P1 = "0b000";
    parameter EXTERNAL_DIVIDE_FACTOR = "0";
    parameter INTFBKDEL_SEL = "DISABLED";
    parameter PMU_WAITFORLOCK = "ENABLED";
    parameter REF_OSC_CTRL = "3P2";
    parameter SIM_FLOAT_PRECISION = "0.0001";
endmodule

module PLLA(INTFBKOP, INTFBKOS, INTFBKOS2, INTFBKOS3, INTFBKOS4, INTFBKOS5, DIR, DIRSEL, LOADREG, DYNROTATE, LMMICLK, LMMIRESET_N, LMMIREQUEST, LMMIWRRD_N, LMMIOFFSET, LMMIWDATA, LMMIRDATA, LMMIRDATAVALID, LMMIREADY, PLLPOWERDOWN_N, REFCK, CLKOP, CLKOS, CLKOS2, CLKOS3, CLKOS4, CLKOS5, ENCLKOP, ENCLKOS, ENCLKOS2, ENCLKOS3, ENCLKOS4, ENCLKOS5, FBKCK, INTLOCK, LEGACY, LEGRDYN, LOCK, PFDDN, PFDUP, PLLRESET, STDBY, REFMUXCK, REGQA, REGQB, REGQB1, CLKOUTDL, ROTDEL, DIRDEL, ROTDELP1, GRAYTEST, BINTEST, DIRDELP1, GRAYACT, BINACT, REFDETRESET, REFDETLOS); //synthesis syn_black_box syn_lib_cell=1
    output INTFBKOP;
    output INTFBKOS;
    output INTFBKOS2;
    output INTFBKOS3;
    output INTFBKOS4;
    output INTFBKOS5;
    input DIR;
    input [2:0] DIRSEL;
    input LOADREG;
    input DYNROTATE;
    input LMMICLK;
    input LMMIRESET_N;
    input LMMIREQUEST;
    input LMMIWRRD_N;
    input [6:0] LMMIOFFSET;
    input [7:0] LMMIWDATA;
    output [7:0] LMMIRDATA;
    output LMMIRDATAVALID;
    output LMMIREADY;
    input PLLPOWERDOWN_N;
    input REFCK;
    output CLKOP;
    output CLKOS;
    output CLKOS2;
    output CLKOS3;
    output CLKOS4;
    output CLKOS5;
    input ENCLKOP;
    input ENCLKOS;
    input ENCLKOS2;
    input ENCLKOS3;
    input ENCLKOS4;
    input ENCLKOS5;
    input FBKCK;
    output INTLOCK;
    input LEGACY;
    output LEGRDYN;
    output LOCK;
    output PFDDN;
    output PFDUP;
    input PLLRESET;
    input STDBY;
    output REFMUXCK;
    output REGQA;
    output REGQB;
    output REGQB1;
    output CLKOUTDL;
    input ROTDEL;
    input DIRDEL;
    input ROTDELP1;
    input [4:0] GRAYTEST;
    input [1:0] BINTEST;
    input DIRDELP1;
    input [4:0] GRAYACT;
    input [1:0] BINACT;
    input REFDETRESET;
    output REFDETLOS;
    parameter BW_CTL_BIAS = "0b0101";
    parameter CLKOP_TRIM = "0b0000";
    parameter CLKOS_TRIM = "0b0000";
    parameter CLKOS2_TRIM = "0b0000";
    parameter CLKOS3_TRIM = "0b0000";
    parameter CLKOS4_TRIM = "0b0000";
    parameter CLKOS5_TRIM = "0b0000";
    parameter CRIPPLE = "5P";
    parameter CSET = "40P";
    parameter DELAY_CTRL = "200PS";
    parameter DELA = "0";
    parameter DELB = "0";
    parameter DELC = "0";
    parameter DELD = "0";
    parameter DELE = "0";
    parameter DELF = "0";
    parameter DIRECTION = "DISABLED";
    parameter DIVA = "0";
    parameter DIVB = "0";
    parameter DIVC = "0";
    parameter DIVD = "0";
    parameter DIVE = "0";
    parameter DIVF = "0";
    parameter DYN_SEL = "0b000";
    parameter DYN_SOURCE = "STATIC";
    parameter ENCLK_CLKOP = "DISABLED";
    parameter ENCLK_CLKOS = "DISABLED";
    parameter ENCLK_CLKOS2 = "DISABLED";
    parameter ENCLK_CLKOS3 = "DISABLED";
    parameter ENCLK_CLKOS4 = "DISABLED";
    parameter ENCLK_CLKOS5 = "DISABLED";
    parameter ENABLE_SYNC = "DISABLED";
    parameter FAST_LOCK_EN = "ENABLED";
    parameter V2I_1V_EN = "DISABLED";
    parameter FBK_CUR_BLE = "0b00000000";
    parameter FBK_EDGE_SEL = "POSITIVE";
    parameter FBK_IF_TIMING_CTL = "0b00";
    parameter FBK_INTEGER_MODE = "DISABLED";
    parameter FBK_MASK = "0b00001000";
    parameter FBK_MMD_DIG = "8";
    parameter FBK_MMD_PULS_CTL = "0b0000";
    parameter FBK_MODE = "0b00";
    parameter FBK_PI_BYPASS = "NOT_BYPASSED";
    parameter FBK_PI_RC = "0b1100";
    parameter FBK_PR_CC = "0b0000";
    parameter FBK_PR_IC = "0b1000";
    parameter FLOAT_CP = "DISABLED";
    parameter FLOCK_CTRL = "2X";
    parameter FLOCK_EN = "ENABLED";
    parameter FLOCK_SRC_SEL = "REFCLK";
    parameter FORCE_FILTER = "DISABLED";
    parameter I_CTRL = "10UA";
    parameter IPI_CMP = "0b1000";
    parameter IPI_CMPN = "0b0011";
    parameter IPI_COMP_EN = "DISABLED";
    parameter IPP_CTRL = "0b1000";
    parameter IPP_SEL = "0b1111";
    parameter KP_VCO = "0b11001";
    parameter LDT_INT_LOCK_STICKY = "DISABLED";
    parameter LDT_LOCK = "1536CYC";
    parameter LDT_LOCK_SEL = "U_FREQ";
    parameter LEGACY_ATT = "DISABLED";
    parameter LOAD_REG = "DISABLED";
    parameter OPENLOOP_EN = "DISABLED";
    parameter PHIA = "0";
    parameter PHIB = "0";
    parameter PHIC = "0";
    parameter PHID = "0";
    parameter PHIE = "0";
    parameter PHIF = "0";
    parameter PLLPDN_EN = "DISABLED";
    parameter PLLPD_N = "UNUSED";
    parameter PLLRESET_ENA = "DISABLED";
    parameter REF_INTEGER_MODE = "DISABLED";
    parameter REF_MASK = "0b00000000";
    parameter REF_MMD_DIG = "8";
    parameter REF_MMD_IN = "0b00001000";
    parameter REF_MMD_PULS_CTL = "0b0000";
    parameter REF_TIMING_CTL = "0b00";
    parameter REFIN_RESET = "SET";
    parameter RESET_LF = "DISABLED";
    parameter ROTATE = "DISABLED";
    parameter SEL_OUTA = "DISABLED";
    parameter SEL_OUTB = "DISABLED";
    parameter SEL_OUTC = "DISABLED";
    parameter SEL_OUTD = "DISABLED";
    parameter SEL_OUTE = "DISABLED";
    parameter SEL_OUTF = "DISABLED";
    parameter SLEEP = "DISABLED";
    parameter SSC_DITHER = "DISABLED";
    parameter SSC_EN_CENTER_IN = "DOWN_TRIANGLE";
    parameter SSC_EN_SDM = "DISABLED";
    parameter SSC_EN_SSC = "DISABLED";
    parameter SSC_F_CODE = "0b000000000000000";
    parameter SSC_N_CODE = "0b000010100";
    parameter SSC_ORDER = "SDM_ORDER2";
    parameter SSC_PI_BYPASS = "NOT_BYPASSED";
    parameter SSC_REG_WEIGHTING_SEL = "0b000";
    parameter SSC_SQUARE_MODE = "DISABLED";
    parameter SSC_STEP_IN = "0b0000000";
    parameter SSC_TBASE = "0b000000000000";
    parameter STDBY_ATT = "DISABLED";
    parameter TRIMOP_BYPASS_N = "BYPASSED";
    parameter TRIMOS_BYPASS_N = "BYPASSED";
    parameter TRIMOS2_BYPASS_N = "BYPASSED";
    parameter TRIMOS3_BYPASS_N = "BYPASSED";
    parameter TRIMOS4_BYPASS_N = "BYPASSED";
    parameter TRIMOS5_BYPASS_N = "BYPASSED";
    parameter V2I_KVCO_SEL = "85";
    parameter V2I_PP_ICTRL = "0b00110";
    parameter V2I_PP_RES = "10K";
    parameter CLKMUX_FB = "CMUX_CLKOP";
    parameter SEL_FBK = "DIVA";
    parameter DIV_DEL = "0b0000001";
    parameter PHASE_SEL_DEL = "0b000";
    parameter PHASE_SEL_DEL_P1 = "0b000";
    parameter EXTERNAL_DIVIDE_FACTOR = "0";
    parameter INTFBKDEL_SEL = "DISABLED";
    parameter PMU_WAITFORLOCK = "ENABLED";
    parameter REF_OSC_CTRL = "3P2";
    parameter REF_COUNTS = "0000";
    parameter SIM_FLOAT_PRECISION = "0.0001";
endmodule

module PREADD9(B, BSIGNED, C, BRS1, BRS2, BLS1, BLS2, BRSS1, BRSS2, BLSS1, BLSS2, PRCASIN, CLK, RSTB, CEB, RSTCL, CECL, BRSO, BLSO, BRSOSGND, BLSOSGND, PRCASOUT, BR, BRSIGNED); //synthesis syn_black_box syn_lib_cell=1
    input [8:0] B;
    input BSIGNED;
    input [9:0] C;
    input [8:0] BRS1;
    input [8:0] BRS2;
    input [8:0] BLS1;
    input [8:0] BLS2;
    input BRSS1;
    input BRSS2;
    input BLSS1;
    input BLSS2;
    input PRCASIN;
    input CLK;
    input RSTB;
    input CEB;
    input RSTCL;
    input CECL;
    output [8:0] BRSO;
    output [8:0] BLSO;
    output BRSOSGND;
    output BLSOSGND;
    output PRCASOUT;
    output [8:0] BR;
    output BRSIGNED;
    parameter SIGNEDSTATIC_EN = "DISABLED";
    parameter SUBSTRACT_EN = "SUBTRACTION";
    parameter CSIGNED = "DISABLED";
    parameter BSIGNED_OPERAND_EN = "DISABLED";
    parameter BYPASS_PREADD9 = "USED";
    parameter REGBYPSBR0 = "REGISTER";
    parameter REGBYPSBR1 = "BYPASS";
    parameter REGBYPSBL = "REGISTER";
    parameter SHIFTBR = "REGISTER";
    parameter SHIFTBL = "REGISTER";
    parameter GSR = "ENABLED";
    parameter PREADDCAS_EN = "DISABLED";
    parameter SR_18BITSHIFT_EN = "DISABLED";
    parameter OPC = "INPUT_B_AS_PREADDER_OPERAND";
    parameter RESET = "SYNC";
endmodule

module PLLREFCS(CLK0, CLK1, SEL, PLLCSOUT); //synthesis syn_black_box syn_lib_cell=1
    input CLK0;
    input CLK1;
    input SEL;
    output PLLCSOUT;
endmodule

module REFMUX(REFCK, ZRSEL3, REFSEL, REFCLK1, REFCLK2); //synthesis syn_black_box syn_lib_cell=1
    output REFCK;
    output ZRSEL3;
    input REFSEL;
    input [7:0] REFCLK1;
    input [7:0] REFCLK2;
    parameter REFSEL_ATT = "MC1";
    parameter SEL1 = "SELECT_REFCLK1";
    parameter SEL_REF2 = "REFCLK2_0";
    parameter SEL_REF1 = "REFCLK1_0";
endmodule

module REG18(PM, PP, CEP, RSTP, CLK); //synthesis syn_black_box syn_lib_cell=1
    input [17:0] PM;
    output [17:0] PP;
    input CEP;
    input RSTP;
    input CLK;
    parameter REGBYPS = "REGISTER";
    parameter GSR = "ENABLED";
    parameter RESET = "SYNC";
endmodule

module SEDC(SEDENABLE, SEDCCOF, SEDCENABLE, SEDCMODE, SEDCSTART, SEDCBUSY, SEDCERR, SEDCERRC, SEDCERRCRC, SEDCERRM, SEDCFRMERRLOC, OSCCLKSEDC, RSTSEDC, SEDCDSRERRLOCCIB); //synthesis syn_black_box syn_lib_cell=1
    input SEDENABLE;
    input SEDCCOF;
    input SEDCENABLE;
    input SEDCMODE;
    input SEDCSTART;
    output SEDCBUSY;
    output SEDCERR;
    output SEDCERRC;
    output SEDCERRCRC;
    output SEDCERRM;
    output [15:0] SEDCFRMERRLOC;
    input OSCCLKSEDC;
    input RSTSEDC;
    output [12:0] SEDCDSRERRLOCCIB;
    parameter SEDCEN = "DIS";
endmodule

module SEIO18(PADDO, DOLP, IOPAD, PADDI, INLP, PADDT, INADC); //synthesis black_box_pad_pin="IOPAD" syn_lib_cell=1
    input PADDO;
    input DOLP;
    inout IOPAD;
    output PADDI;
    output INLP;
    input PADDT;
    output INADC;
    parameter PULLMODE = "DOWN";
    parameter MIPI = "DISABLED";
    parameter ENADC_IN = "DISABLED";
endmodule

module SEIO33(IOPAD, PADDI, PADDO, PADDT, I3CRESEN, I3CWKPU); //synthesis black_box_pad_pin="IOPAD" syn_lib_cell=1
    inout IOPAD;
    output PADDI;
    input PADDO;
    input PADDT;
    input I3CRESEN;
    input I3CWKPU;
    parameter PULLMODE = "DOWN";
endmodule

module SGMIICDR(LMMICLK, LMMIRESET_N, LMMIREQUEST, LMMIWRRD_N, LMMIOFFSET, LMMIWDATA, LMMIRDATA, LMMIRDATAVALID, LMMIREADY, DCALIRST, DFACQRST, RRST, SPCLK, SRCLK, SRXD, RSTBFBW, RSTBRXF, SGMIIIN, SREFCLK, CDRLOL); //synthesis syn_black_box syn_lib_cell=1
    input LMMICLK;
    input LMMIRESET_N;
    input LMMIREQUEST;
    input LMMIWRRD_N;
    input [3:0] LMMIOFFSET;
    input [7:0] LMMIWDATA;
    output [7:0] LMMIRDATA;
    output LMMIRDATAVALID;
    output LMMIREADY;
    input DCALIRST;
    input DFACQRST;
    input RRST;
    input SPCLK;
    output SRCLK;
    output [9:0] SRXD;
    input RSTBFBW;
    input RSTBRXF;
    input SGMIIIN;
    input SREFCLK;
    output CDRLOL;
    parameter GSR = "ENABLED";
    parameter DCOITUNE4LSB = "0_PERCENT";
    parameter DCOCTLGI = "60_PERCENT";
    parameter DCOSTEP = "17_PERCENT";
    parameter DCOCALDIV = "100_PERCENT";
    parameter DCOIOSTUNE = "49_PERCENT";
    parameter DCOFLTDAC = "181MHZ";
    parameter DCOSTARTVAL = "100_PERCENT";
    parameter DCONUOFLSB = "60_PERCENT";
    parameter RPWDNB = "POWER_UP";
    parameter CDR_CNT4SEL = "BY_4";
    parameter DCOITUNE = "100_PERCENT";
    parameter BAND_THRESHOLD = "0b000000";
    parameter AUTO_FACQ_EN = "ENABLED";
    parameter AUTO_CALIB_EN = "ENABLED";
    parameter CDR_LOL_SET = "2000_PPM";
    parameter FC2DCO_FLOOP = "DISABLED";
    parameter FC2DCO_DLOOP = "DISABLED";
    parameter CALIB_TIME_SEL = "24_CYC";
    parameter CALIB_CK_MODE = "BY_2";
    parameter BAND_CALIB_MODE = "256_FDBK_CLK_CYC";
    parameter REG_BAND_SEL = "0b10101";
    parameter REG_BAND_OFFSET = "0b0000";
    parameter REG_IDAC_SEL = "0b10000000";
    parameter LB_CTL = "DISABLED";
    parameter REG_IDAC_EN = "DISABLED";
    parameter ATDCFG = "0_PS";
    parameter ATDDLY = "0_PS";
    parameter BDAVOID_ENB = "ENABLED";
    parameter BYPASSATD = "NOT_BYPASS";
    parameter DCOIUPDNX2 = "2X";
    parameter IDAC_EN = "DISABLED";
    parameter FB_CLK_DIV = "0b010";
    parameter EN_RECALIB = "ENABLED";
endmodule

module SP16K_MODE(DI0, DI1, DI2, DI3, DI4, DI5, DI6, DI7, DI8, DI9, DI10, DI11, DI12, DI13, DI14, DI15, DI16, DI17, AD0, AD1, AD2, AD3, AD4, AD5, AD6, AD7, AD8, AD9, AD10, AD11, AD12, AD13, CLK, CE, WE, CS0, CS1, CS2, RST, DO0, DO1, DO2, DO3, DO4, DO5, DO6, DO7, DO8, DO9, DO10, DO11, DO12, DO13, DO14, DO15, DO16, DO17); //synthesis syn_black_box syn_lib_cell=1
    input DI0;
    input DI1;
    input DI2;
    input DI3;
    input DI4;
    input DI5;
    input DI6;
    input DI7;
    input DI8;
    input DI9;
    input DI10;
    input DI11;
    input DI12;
    input DI13;
    input DI14;
    input DI15;
    input DI16;
    input DI17;
    input AD0;
    input AD1;
    input AD2;
    input AD3;
    input AD4;
    input AD5;
    input AD6;
    input AD7;
    input AD8;
    input AD9;
    input AD10;
    input AD11;
    input AD12;
    input AD13;
    input CLK;
    input CE;
    input WE;
    input CS0;
    input CS1;
    input CS2;
    input RST;
    output DO0;
    output DO1;
    output DO2;
    output DO3;
    output DO4;
    output DO5;
    output DO6;
    output DO7;
    output DO8;
    output DO9;
    output DO10;
    output DO11;
    output DO12;
    output DO13;
    output DO14;
    output DO15;
    output DO16;
    output DO17;
    parameter DATA_WIDTH = "X18";
    parameter OUTREG = "BYPASSED";
    parameter RESETMODE = "SYNC";
    parameter GSR = "ENABLED";
    parameter INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter CSDECODE = "000";
    parameter ASYNC_RST_RELEASE = "SYNC";
    parameter INIT_DATA = "STATIC";
endmodule

module SP16K(DI, AD, CLK, CE, WE, CS, RST, DO); //synthesis syn_black_box syn_lib_cell=1
    input [17:0] DI;
    input [13:0] AD;
    input CLK;
    input CE;
    input WE;
    input [2:0] CS;
    input RST;
    output [17:0] DO;
    parameter DATA_WIDTH = "X18";
    parameter OUTREG = "BYPASSED";
    parameter RESETMODE = "SYNC";
    parameter GSR = "ENABLED";
    parameter INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter CSDECODE = "000";
    parameter ASYNC_RST_RELEASE = "SYNC";
    parameter INIT_DATA = "STATIC";
endmodule

module SP512K(DI, AD, CLK, CE, WE, CS, RSTOUT, CEOUT, BYTEEN_N, DO, ERRDECA, ERRDECB); //synthesis syn_black_box syn_lib_cell=1
    input [31:0] DI;
    input [13:0] AD;
    input CLK;
    input CE;
    input WE;
    input CS;
    input RSTOUT;
    input CEOUT;
    input [3:0] BYTEEN_N;
    output [31:0] DO;
    output [1:0] ERRDECA;
    output [1:0] ERRDECB;
    parameter OUTREG = "NO_REG";
    parameter GSR = "ENABLED";
    parameter RESETMODE = "SYNC";
    parameter INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_40 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_41 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_42 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_43 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_44 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_45 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_46 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_47 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_48 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_49 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_4A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_4B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_4C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_4D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_4E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_4F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_50 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_51 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_52 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_53 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_54 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_55 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_56 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_57 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_58 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_59 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_5A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_5B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_5C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_5D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_5E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_5F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_60 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_61 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_62 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_63 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_64 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_65 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_66 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_67 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_68 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_69 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_6A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_6B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_6C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_6D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_6E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_6F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_70 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_71 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_72 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_73 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_74 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_75 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_76 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_77 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_78 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_79 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_7A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_7B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_7C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_7D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_7E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter INITVAL_7F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    parameter ASYNC_RESET_RELEASE = "SYNC";
    parameter ECC_BYTE_SEL = "ECC_EN";
endmodule

module TSHX2DQS(T0, T1, DQSW, ECLK, SCLK, RST, Q); //synthesis syn_black_box syn_lib_cell=1
    input T0;
    input T1;
    input DQSW;
    input ECLK;
    input SCLK;
    input RST;
    output Q;
    parameter GSR = "ENABLED";
endmodule

module TSHX2DQ(T0, T1, DQSW270, ECLK, SCLK, RST, Q); //synthesis syn_black_box syn_lib_cell=1
    input T0;
    input T1;
    input DQSW270;
    input ECLK;
    input SCLK;
    input RST;
    output Q;
    parameter GSR = "ENABLED";
endmodule

module TSHX4DQS(T0, T1, T2, T3, DQSW, ECLK, SCLK, RST, Q); //synthesis syn_black_box syn_lib_cell=1
    input T0;
    input T1;
    input T2;
    input T3;
    input DQSW;
    input ECLK;
    input SCLK;
    input RST;
    output Q;
    parameter GSR = "ENABLED";
endmodule

module TSHX4DQ(T0, T1, T2, T3, DQSW270, ECLK, SCLK, RST, Q); //synthesis syn_black_box syn_lib_cell=1
    input T0;
    input T1;
    input T2;
    input T3;
    input DQSW270;
    input ECLK;
    input SCLK;
    input RST;
    output Q;
    parameter GSR = "ENABLED";
endmodule

module WDT(WDTRELOAD, WDT_CLK, WDT_RST); //synthesis syn_noprune=1 syn_lib_cell=1
    input WDTRELOAD;
    input WDT_CLK;
    input WDT_RST;
    parameter WDTEN = "DIS";
    parameter WDTMODE = "SINGLE";
    parameter WDTVALUE = "0b000000000000000000";
endmodule

module MIPI(AP, AN, TP, TN, HSRXEN, HSTXEN, BP, BN, OLSP, OLSN, OHS, IHS); //synthesis syn_black_box black_box_pad_pin="BP,BN" syn_lib_cell=1
    inout BP;
    inout BN;
    input AP;
    input AN;
    input TP;
    input TN;
    input IHS;
    input HSRXEN;
    input HSTXEN;
    output OHS;
    output OLSP;
    output OLSN;
    parameter MIPI_ID = "0";
endmodule


module CONFIG_IP_CORE (
CFGDONECIB, CIBTSALL, FREEZEIOCIB, LASTADDRCIB15, LASTADDRCIB14, LASTADDRCIB13,
LASTADDRCIB12, LASTADDRCIB11, LASTADDRCIB10, LASTADDRCIB9, LASTADDRCIB8,
LASTADDRCIB7, LASTADDRCIB6, LASTADDRCIB5, LASTADDRCIB4, LASTADDRCIB3, LASTADDRCIB2,
LASTADDRCIB1, LASTADDRCIB0, MBISTENABLEN, MBISTRRMATCH, MBISTTRRAEN) ;  //synthesis  syn_black_box  syn_lib_cell=1

        output CFGDONECIB;
        input CIBTSALL;
        output FREEZEIOCIB;
        output LASTADDRCIB15;
        output LASTADDRCIB14;
        output LASTADDRCIB13;
        output LASTADDRCIB12;
        output LASTADDRCIB11;
        output LASTADDRCIB10;
        output LASTADDRCIB9;
        output LASTADDRCIB8;
        output LASTADDRCIB7;
        output LASTADDRCIB6;
        output LASTADDRCIB5;
        output LASTADDRCIB4;
        output LASTADDRCIB3;
        output LASTADDRCIB2;
        output LASTADDRCIB1;
        output LASTADDRCIB0;
        input MBISTENABLEN;
        output MBISTRRMATCH;
        input MBISTTRRAEN;

        parameter DONEPHASE = "DIS";
        parameter DSRFCTRL = "0b00";
        parameter ENTSALL = "DIS";
        parameter MCCFGUSEREN = "DIS";
        parameter MCCIBINT = "DIS";
        parameter MCHSEUSEREN = "DIS";
        parameter MCJTAGDISABLE = "EN";
        parameter MCPERSISTUI2C = "DIS";
        parameter MCSPARE = "0b00000";
        parameter MCUCLKSEL = "DIS";
        parameter MCUI2CAFWKUP = "DIS";
        parameter PERSISTI2C = "DIS";
        parameter PERSISTI3C = "DIS";
        parameter PERSISTMQUAD = "DIS";
        parameter PERSISTMSPI = "DIS";
        parameter PERSISTSHEXA = "DIS";
        parameter PERSISTSOCTA = "DIS";
        parameter PERSISTSQUAD = "DIS";
        parameter PERSISTSSPI = "DIS";
        parameter PERSISTWKUP = "DIS";
        parameter PPTQOUT = "0b0000";
        parameter SCANEN = "DIS";
        parameter SYNCEXTDONE = "DIS";
        parameter TRANECI = "DIS";
        parameter TRANHSE = "DIS";
        parameter TRANSBI = "DIS";
        parameter TSALLINV = "NINV";
        parameter WLSLEW = "DIS";

endmodule



module TSALLA(TSALL); //synthesis syn_black_box syn_noprune=1 syn_lib_cell=1
    input TSALL;
endmodule



module OSCA(HFOUTEN, HFSDSCEN, HFCLKOUT, LFCLKOUT, HFCLKCFG, HFSDCOUT); //synthesis syn_black_box syn_lib_cell=1

    input HFOUTEN;
    input HFSDSCEN;
    output HFCLKOUT;
    output LFCLKOUT;
    output HFCLKCFG;
    output HFSDCOUT;

    parameter HF_CLK_DIV = "1";
    parameter HF_SED_SEC_DIV = "1";
    parameter HF_OSC_EN = "ENABLED";
    parameter LF_OUTPUT_EN = "DISABLED";
endmodule




module OSC(HFCLKOUT, HFSDSCEN, LFCLKOUT, HFSDCOUT, HSE_CLK, JTAG_LRST_N, LMMI_CLK, LMMI_CLK_O, LMMI_LRST_N, LMMI_RST, SEDC_CLK, SEDC_LRST_N, SEDC_RST, CFG_CLK, SMCLK_RST, WDT_CLK, WDT_LRST_N, WDT_RST); //synthesis syn_black_box syn_lib_cell=1
    output HFCLKOUT;
    input HFSDSCEN;
    output LFCLKOUT;
    output HFSDCOUT;
	output HSE_CLK;
	input JTAG_LRST_N;
	input LMMI_CLK;
	output LMMI_CLK_O;
	input LMMI_LRST_N;
	output LMMI_RST;
	input SEDC_CLK;
	input SEDC_LRST_N;
	output SEDC_RST;
	output CFG_CLK;
	output SMCLK_RST;
	output WDT_CLK;
	input WDT_LRST_N;
	output WDT_RST;
    parameter DTR_EN = "ENABLED";
    parameter HF_CLK_DIV = "1";
    parameter HF_SED_SEC_DIV = "1";
    parameter HF_FABRIC_EN = "DISABLED";
    parameter HF_OSC_EN = "ENABLED";
    parameter HFDIV_FABRIC_EN = "ENABLED";
    parameter LF_FABRIC_EN = "DISABLED";
    parameter LF_OUTPUT_EN = "DISABLED";
    parameter DEBUG_N = "DISABLED";
	parameter MCJTAGGSRNDIS = "EN";
	parameter MCLMMIGSRNDIS = "EN";
	parameter MCSEDCGSRNDIS = "EN";
	parameter MCWDTGSRNDIS = "EN";
	parameter SMCLK_DIV = "3";
endmodule

module ACC54_CORE (SFTCTRL3, SFTCTRL2, SFTCTRL1, SFTCTRL0, DSPIN53, DSPIN52, DSPIN51, DSPIN50, DSPIN49, DSPIN48, DSPIN47, DSPIN46, DSPIN45, DSPIN44, DSPIN43, DSPIN42, DSPIN41, DSPIN40, DSPIN39, DSPIN38, DSPIN37, DSPIN36, DSPIN35, DSPIN34, DSPIN33, DSPIN32, DSPIN31, DSPIN30, DSPIN29, DSPIN28, DSPIN27, DSPIN26, DSPIN25, DSPIN24, DSPIN23, DSPIN22, DSPIN21, DSPIN20, DSPIN19, DSPIN18, DSPIN17, DSPIN16, DSPIN15, DSPIN14, DSPIN13, DSPIN12, DSPIN11, DSPIN10, DSPIN9, DSPIN8, DSPIN7, DSPIN6, DSPIN5, DSPIN4, DSPIN3, DSPIN2, DSPIN1, DSPIN0, PP71, PP70, PP69, PP68, PP67, PP66, PP65, PP64, PP63, PP62, PP61, PP60, PP59, PP58, PP57, PP56, PP55, PP54, PP53, PP52, PP51, PP50, PP49, PP48, PP47, PP46, PP45, PP44, PP43, PP42, PP41, PP40, PP39, PP38, PP37, PP36, PP35, PP34, PP33, PP32, PP31, PP30, PP29, PP28, PP27, PP26, PP25, PP24, PP23, PP22, PP21, PP20, PP19, PP18, PP17, PP16, PP15, PP14, PP13, PP12, PP11, PP10, PP9, PP8, PP7, PP6, PP5, PP4, PP3, PP2, PP1, PP0, CINPUT53, CINPUT52, CINPUT51, CINPUT50, CINPUT49, CINPUT48, CINPUT47, CINPUT46, CINPUT45, CINPUT44, CINPUT43, CINPUT42, CINPUT41, CINPUT40, CINPUT39, CINPUT38, CINPUT37, CINPUT36, CINPUT35, CINPUT34, CINPUT33, CINPUT32, CINPUT31, CINPUT30, CINPUT29, CINPUT28, CINPUT27, CINPUT26, CINPUT25, CINPUT24, CINPUT23, CINPUT22, CINPUT21, CINPUT20, CINPUT19, CINPUT18, CINPUT17, CINPUT16, CINPUT15, CINPUT14, CINPUT13, CINPUT12, CINPUT11, CINPUT10, CINPUT9, CINPUT8, CINPUT7, CINPUT6, CINPUT5, CINPUT4, CINPUT3, CINPUT2, CINPUT1, CINPUT0, LOAD, M9ADDSUB1, M9ADDSUB0, ADDSUB1, ADDSUB0, CIN, CASIN1, CASIN0, CEO, RSTO, CEC, RSTC, CLK, SIGNEDI, SUM135, SUM134, SUM133, SUM132, SUM131, SUM130, SUM129, SUM128, SUM127, SUM126, SUM125, SUM124, SUM123, SUM122, SUM121, SUM120, SUM119, SUM118, SUM117, SUM116, SUM115, SUM114, SUM113, SUM112, SUM111, SUM110, SUM19, SUM18, SUM17, SUM16, SUM15, SUM14, SUM13, SUM12, SUM11, SUM10, SUM035, SUM034, SUM033, SUM032, SUM031, SUM030, SUM029, SUM028, SUM027, SUM026, SUM025, SUM024, SUM023, SUM022, SUM021, SUM020, SUM019, SUM018, SUM017, SUM016, SUM015, SUM014, SUM013, SUM012, SUM011, SUM010, SUM09, SUM08, SUM07, SUM06, SUM05, SUM04, SUM03, SUM02, SUM01, SUM00, DSPOUT53, DSPOUT52, DSPOUT51, DSPOUT50, DSPOUT49, DSPOUT48, DSPOUT47, DSPOUT46, DSPOUT45, DSPOUT44, DSPOUT43, DSPOUT42, DSPOUT41, DSPOUT40, DSPOUT39, DSPOUT38, DSPOUT37, DSPOUT36, DSPOUT35, DSPOUT34, DSPOUT33, DSPOUT32, DSPOUT31, DSPOUT30, DSPOUT29, DSPOUT28, DSPOUT27, DSPOUT26, DSPOUT25, DSPOUT24, DSPOUT23, DSPOUT22, DSPOUT21, DSPOUT20, DSPOUT19, DSPOUT18, DSPOUT17, DSPOUT16, DSPOUT15, DSPOUT14, DSPOUT13, DSPOUT12, DSPOUT11, DSPOUT10, DSPOUT9, DSPOUT8, DSPOUT7, DSPOUT6, DSPOUT5, DSPOUT4, DSPOUT3, DSPOUT2, DSPOUT1, DSPOUT0, CASCOUT1, CASCOUT0, ROUNDEN, CECIN, CECTRL, RSTCIN, RSTCTRL); //synthesis syn_black_box syn_lib_cell=1

	input SFTCTRL3;
	input SFTCTRL2;
	input SFTCTRL1;
	input SFTCTRL0;
	input DSPIN53;
	input DSPIN52;
	input DSPIN51;
	input DSPIN50;
	input DSPIN49;
	input DSPIN48;
	input DSPIN47;
	input DSPIN46;
	input DSPIN45;
	input DSPIN44;
	input DSPIN43;
	input DSPIN42;
	input DSPIN41;
	input DSPIN40;
	input DSPIN39;
	input DSPIN38;
	input DSPIN37;
	input DSPIN36;
	input DSPIN35;
	input DSPIN34;
	input DSPIN33;
	input DSPIN32;
	input DSPIN31;
	input DSPIN30;
	input DSPIN29;
	input DSPIN28;
	input DSPIN27;
	input DSPIN26;
	input DSPIN25;
	input DSPIN24;
	input DSPIN23;
	input DSPIN22;
	input DSPIN21;
	input DSPIN20;
	input DSPIN19;
	input DSPIN18;
	input DSPIN17;
	input DSPIN16;
	input DSPIN15;
	input DSPIN14;
	input DSPIN13;
	input DSPIN12;
	input DSPIN11;
	input DSPIN10;
	input DSPIN9;
	input DSPIN8;
	input DSPIN7;
	input DSPIN6;
	input DSPIN5;
	input DSPIN4;
	input DSPIN3;
	input DSPIN2;
	input DSPIN1;
	input DSPIN0;
	input PP71;
	input PP70;
	input PP69;
	input PP68;
	input PP67;
	input PP66;
	input PP65;
	input PP64;
	input PP63;
	input PP62;
	input PP61;
	input PP60;
	input PP59;
	input PP58;
	input PP57;
	input PP56;
	input PP55;
	input PP54;
	input PP53;
	input PP52;
	input PP51;
	input PP50;
	input PP49;
	input PP48;
	input PP47;
	input PP46;
	input PP45;
	input PP44;
	input PP43;
	input PP42;
	input PP41;
	input PP40;
	input PP39;
	input PP38;
	input PP37;
	input PP36;
	input PP35;
	input PP34;
	input PP33;
	input PP32;
	input PP31;
	input PP30;
	input PP29;
	input PP28;
	input PP27;
	input PP26;
	input PP25;
	input PP24;
	input PP23;
	input PP22;
	input PP21;
	input PP20;
	input PP19;
	input PP18;
	input PP17;
	input PP16;
	input PP15;
	input PP14;
	input PP13;
	input PP12;
	input PP11;
	input PP10;
	input PP9;
	input PP8;
	input PP7;
	input PP6;
	input PP5;
	input PP4;
	input PP3;
	input PP2;
	input PP1;
	input PP0;
	input CINPUT53;
	input CINPUT52;
	input CINPUT51;
	input CINPUT50;
	input CINPUT49;
	input CINPUT48;
	input CINPUT47;
	input CINPUT46;
	input CINPUT45;
	input CINPUT44;
	input CINPUT43;
	input CINPUT42;
	input CINPUT41;
	input CINPUT40;
	input CINPUT39;
	input CINPUT38;
	input CINPUT37;
	input CINPUT36;
	input CINPUT35;
	input CINPUT34;
	input CINPUT33;
	input CINPUT32;
	input CINPUT31;
	input CINPUT30;
	input CINPUT29;
	input CINPUT28;
	input CINPUT27;
	input CINPUT26;
	input CINPUT25;
	input CINPUT24;
	input CINPUT23;
	input CINPUT22;
	input CINPUT21;
	input CINPUT20;
	input CINPUT19;
	input CINPUT18;
	input CINPUT17;
	input CINPUT16;
	input CINPUT15;
	input CINPUT14;
	input CINPUT13;
	input CINPUT12;
	input CINPUT11;
	input CINPUT10;
	input CINPUT9;
	input CINPUT8;
	input CINPUT7;
	input CINPUT6;
	input CINPUT5;
	input CINPUT4;
	input CINPUT3;
	input CINPUT2;
	input CINPUT1;
	input CINPUT0;
	input LOAD;
	input M9ADDSUB1;
	input M9ADDSUB0;
	input ADDSUB1;
	input ADDSUB0;
	input CIN;
	input CASIN1;
	input CASIN0;
	input CEO;
	input RSTO;
	input CEC;
	input RSTC;
	input CLK;
	input SIGNEDI;
	output SUM135;
	output SUM134;
	output SUM133;
	output SUM132;
	output SUM131;
	output SUM130;
	output SUM129;
	output SUM128;
	output SUM127;
	output SUM126;
	output SUM125;
	output SUM124;
	output SUM123;
	output SUM122;
	output SUM121;
	output SUM120;
	output SUM119;
	output SUM118;
	output SUM117;
	output SUM116;
	output SUM115;
	output SUM114;
	output SUM113;
	output SUM112;
	output SUM111;
	output SUM110;
	output SUM19;
	output SUM18;
	output SUM17;
	output SUM16;
	output SUM15;
	output SUM14;
	output SUM13;
	output SUM12;
	output SUM11;
	output SUM10;
	output SUM035;
	output SUM034;
	output SUM033;
	output SUM032;
	output SUM031;
	output SUM030;
	output SUM029;
	output SUM028;
	output SUM027;
	output SUM026;
	output SUM025;
	output SUM024;
	output SUM023;
	output SUM022;
	output SUM021;
	output SUM020;
	output SUM019;
	output SUM018;
	output SUM017;
	output SUM016;
	output SUM015;
	output SUM014;
	output SUM013;
	output SUM012;
	output SUM011;
	output SUM010;
	output SUM09;
	output SUM08;
	output SUM07;
	output SUM06;
	output SUM05;
	output SUM04;
	output SUM03;
	output SUM02;
	output SUM01;
	output SUM00;
	output DSPOUT53;
	output DSPOUT52;
	output DSPOUT51;
	output DSPOUT50;
	output DSPOUT49;
	output DSPOUT48;
	output DSPOUT47;
	output DSPOUT46;
	output DSPOUT45;
	output DSPOUT44;
	output DSPOUT43;
	output DSPOUT42;
	output DSPOUT41;
	output DSPOUT40;
	output DSPOUT39;
	output DSPOUT38;
	output DSPOUT37;
	output DSPOUT36;
	output DSPOUT35;
	output DSPOUT34;
	output DSPOUT33;
	output DSPOUT32;
	output DSPOUT31;
	output DSPOUT30;
	output DSPOUT29;
	output DSPOUT28;
	output DSPOUT27;
	output DSPOUT26;
	output DSPOUT25;
	output DSPOUT24;
	output DSPOUT23;
	output DSPOUT22;
	output DSPOUT21;
	output DSPOUT20;
	output DSPOUT19;
	output DSPOUT18;
	output DSPOUT17;
	output DSPOUT16;
	output DSPOUT15;
	output DSPOUT14;
	output DSPOUT13;
	output DSPOUT12;
	output DSPOUT11;
	output DSPOUT10;
	output DSPOUT9;
	output DSPOUT8;
	output DSPOUT7;
	output DSPOUT6;
	output DSPOUT5;
	output DSPOUT4;
	output DSPOUT3;
	output DSPOUT2;
	output DSPOUT1;
	output DSPOUT0;
	output CASCOUT1;
	output CASCOUT0;
	input ROUNDEN;
	input CECIN;
	input CECTRL;
	input RSTCIN;
	input RSTCTRL;

	parameter SIGN = "DISABLED";
	parameter M9ADDSUB_CTRL = "ADDITION";
	parameter ADDSUB_CTRL = "ADD_ADD_CTRL_54_BIT_ADDER";
	parameter STATICOPCODE_EN = "DISABLED";
	parameter OUTREGBYPS = "REGISTER";
	parameter GSR = "ENABLED";
	parameter PROGCONST = "0b000000000000000000000000000000000000000000000000000000";
	parameter CONSTSEL = "BYPASS";
	parameter DSPCASCADE = "DISABLED";
	parameter ACC108CASCADE = "BYPASSCASCADE";
	parameter ACCUMODE = "MODE0";
	parameter ACCUBYPS = "USED";
	parameter CREGBYPS1 = "REGISTER";
	parameter CREGBYPS2 = "REGISTER";
	parameter CREGBYPS3 = "REGISTER";
	parameter CINREGBYPS1 = "REGISTER";
	parameter CINREGBYPS2 = "REGISTER";
	parameter CINREGBYPS3 = "REGISTER";
	parameter LOADREGBYPS1 = "REGISTER";
	parameter LOADREGBYPS2 = "REGISTER";
	parameter LOADREGBYPS3 = "REGISTER";
	parameter M9ADDSUBREGBYPS1 = "REGISTER";
	parameter M9ADDSUBREGBYPS2 = "REGISTER";
	parameter M9ADDSUBREGBYPS3 = "REGISTER";
	parameter ADDSUBSIGNREGBYPS1 = "REGISTER";
	parameter ADDSUBSIGNREGBYPS2 = "REGISTER";
	parameter ADDSUBSIGNREGBYPS3 = "REGISTER";
	parameter ROUNDHALFUP = "DISABLED";
	parameter ROUNDRTZI = "ROUND_TO_ZERO";
	parameter ROUNDBIT = "ROUND_TO_BIT0";
	parameter CASCOUTREGBYPS = "REGISTER";
	parameter SFTEN = "DISABLED";
	parameter RESET = "SYNC";

endmodule

module ADC_CORE (ADCEN, CAL, CALRDY, CHAEN, CHASEL3, CHASEL2, CHASEL1, CHASEL0, CHBEN, CHBSEL3, CHBSEL2, CHBSEL1, CHBSEL0, CLKDCLK, CLKFAB, COG, COMP1IN, COMP1IP, COMP1OL, COMP2IN, COMP2IP, COMP2OL, COMP3IN, COMP3IP, COMP3OL, CONVSTOP, DA11, DA10, DA9, DA8, DA7, DA6, DA5, DA4, DA3, DA2, DA1, DA0, DB11, DB10, DB9, DB8, DB7, DB6, DB5, DB4, DB3, DB2, DB1, DB0, DN1, DN0, DP1, DP0, EOC, GPION15, GPION14, GPION13, GPION12, GPION11, GPION10, GPION9, GPION8, GPION7, GPION6, GPION5, GPION4, GPION3, GPION2, GPION1, GPION0, GPIOP15, GPIOP14, GPIOP13, GPIOP12, GPIOP11, GPIOP10, GPIOP9, GPIOP8, GPIOP7, GPIOP6, GPIOP5, GPIOP4, GPIOP3, GPIOP2, GPIOP1, GPIOP0, RESETN, RSTN, RSVDH, RSVDL, SOC, COMP1O, COMP2O, COMP3O); //synthesis syn_black_box black_box_pad_pin="DN1,DN0,DP1,DP0" syn_lib_cell=1

	input ADCEN;
	input CAL;
	output CALRDY;
	input CHAEN;
	input CHASEL3;
	input CHASEL2;
	input CHASEL1;
	input CHASEL0;
	input CHBEN;
	input CHBSEL3;
	input CHBSEL2;
	input CHBSEL1;
	input CHBSEL0;
	input CLKDCLK;
	input CLKFAB;
	output COG;
	input COMP1IN;
	input COMP1IP;
	output COMP1OL;
	input COMP2IN;
	input COMP2IP;
	output COMP2OL;
	input COMP3IN;
	input COMP3IP;
	output COMP3OL;
	input CONVSTOP;
	output DA11;
	output DA10;
	output DA9;
	output DA8;
	output DA7;
	output DA6;
	output DA5;
	output DA4;
	output DA3;
	output DA2;
	output DA1;
	output DA0;
	output DB11;
	output DB10;
	output DB9;
	output DB8;
	output DB7;
	output DB6;
	output DB5;
	output DB4;
	output DB3;
	output DB2;
	output DB1;
	output DB0;
	input DN1;
	input DN0;
	input DP1;
	input DP0;
	output EOC;
	input GPION15;
	input GPION14;
	input GPION13;
	input GPION12;
	input GPION11;
	input GPION10;
	input GPION9;
	input GPION8;
	input GPION7;
	input GPION6;
	input GPION5;
	input GPION4;
	input GPION3;
	input GPION2;
	input GPION1;
	input GPION0;
	input GPIOP15;
	input GPIOP14;
	input GPIOP13;
	input GPIOP12;
	input GPIOP11;
	input GPIOP10;
	input GPIOP9;
	input GPIOP8;
	input GPIOP7;
	input GPIOP6;
	input GPIOP5;
	input GPIOP4;
	input GPIOP3;
	input GPIOP2;
	input GPIOP1;
	input GPIOP0;
	input RESETN;
	input RSTN;
	input RSVDH;
	input RSVDL;
	input SOC;
	output COMP1O;
	output COMP2O;
	output COMP3O;

	parameter ADC_ENP = "ENABLED";
	parameter CLK_DIV = "2";
	parameter CTLCOMPSW1 = "DISABLED";
	parameter CTLCOMPSW2 = "DISABLED";
	parameter CTLCOMPSW3 = "DISABLED";
	parameter DF = "STRAIGHT_BINARY";
	parameter EN_COMP1 = "ENABLED";
	parameter EN_COMP2 = "ENABLED";
	parameter EN_COMP3 = "ENABLED";
	parameter OMA = "BIPOLAR";
	parameter OMB = "BIPOLAR";
	parameter REFBUFAEN = "ENABLED";
	parameter REFBUFBEN = "ENABLED";
	parameter SLEEP = "DISABLED";
	parameter VREFACFG = "1P0_TO_1P2";
	parameter VREFASEL = "INTERNAL";
	parameter VREFBCFG = "1P0_TO_1P2";
	parameter VREFBSEL = "INTERNAL";

endmodule

module ALUREG_CORE (OPCGLOADCLK, ALUCLK, ALUFLAGC, ALUFLAGV, ALUFLAGZ, ALUFORWARDA, ALUFORWARDB, ALUIREGEN, ALUOREGEN, ALURST, DATAA31, DATAA30, DATAA29, DATAA28, DATAA27, DATAA26, DATAA25, DATAA24, DATAA23, DATAA22, DATAA21, DATAA20, DATAA19, DATAA18, DATAA17, DATAA16, DATAA15, DATAA14, DATAA13, DATAA12, DATAA11, DATAA10, DATAA9, DATAA8, DATAA7, DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0, DATAB31, DATAB30, DATAB29, DATAB28, DATAB27, DATAB26, DATAB25, DATAB24, DATAB23, DATAB22, DATAB21, DATAB20, DATAB19, DATAB18, DATAB17, DATAB16, DATAB15, DATAB14, DATAB13, DATAB12, DATAB11, DATAB10, DATAB9, DATAB8, DATAB7, DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0, DATAC4, DATAC3, DATAC2, DATAC1, DATAC0, OPC6, OPC5, OPC4, OPC3, OPC2, OPC1, OPC0, OPCCUSTOM, RADDRA4, RADDRA3, RADDRA2, RADDRA1, RADDRA0, RADDRB4, RADDRB3, RADDRB2, RADDRB1, RADDRB0, RDATAA31, RDATAA30, RDATAA29, RDATAA28, RDATAA27, RDATAA26, RDATAA25, RDATAA24, RDATAA23, RDATAA22, RDATAA21, RDATAA20, RDATAA19, RDATAA18, RDATAA17, RDATAA16, RDATAA15, RDATAA14, RDATAA13, RDATAA12, RDATAA11, RDATAA10, RDATAA9, RDATAA8, RDATAA7, RDATAA6, RDATAA5, RDATAA4, RDATAA3, RDATAA2, RDATAA1, RDATAA0, RDATAB31, RDATAB30, RDATAB29, RDATAB28, RDATAB27, RDATAB26, RDATAB25, RDATAB24, RDATAB23, RDATAB22, RDATAB21, RDATAB20, RDATAB19, RDATAB18, RDATAB17, RDATAB16, RDATAB15, RDATAB14, RDATAB13, RDATAB12, RDATAB11, RDATAB10, RDATAB9, RDATAB8, RDATAB7, RDATAB6, RDATAB5, RDATAB4, RDATAB3, RDATAB2, RDATAB1, RDATAB0, REGCLK, REGCLKEN, REGRST, RESULT31, RESULT30, RESULT29, RESULT28, RESULT27, RESULT26, RESULT25, RESULT24, RESULT23, RESULT22, RESULT21, RESULT20, RESULT19, RESULT18, RESULT17, RESULT16, RESULT15, RESULT14, RESULT13, RESULT12, RESULT11, RESULT10, RESULT9, RESULT8, RESULT7, RESULT6, RESULT5, RESULT4, RESULT3, RESULT2, RESULT1, RESULT0, SCANCLK, SCANRST, WADDR4, WADDR3, WADDR2, WADDR1, WADDR0, WDROTATE1, WDROTATE0, WDSIGNEXT, WDSIZE1, WDSIZE0, WDATA31, WDATA30, WDATA29, WDATA28, WDATA27, WDATA26, WDATA25, WDATA24, WDATA23, WDATA22, WDATA21, WDATA20, WDATA19, WDATA18, WDATA17, WDATA16, WDATA15, WDATA14, WDATA13, WDATA12, WDATA11, WDATA10, WDATA9, WDATA8, WDATA7, WDATA6, WDATA5, WDATA4, WDATA3, WDATA2, WDATA1, WDATA0, WREN); //synthesis syn_black_box syn_lib_cell=1

	input OPCGLOADCLK;
	input ALUCLK;
	output ALUFLAGC;
	output ALUFLAGV;
	output ALUFLAGZ;
	input ALUFORWARDA;
	input ALUFORWARDB;
	input ALUIREGEN;
	input ALUOREGEN;
	input ALURST;
	input DATAA31;
	input DATAA30;
	input DATAA29;
	input DATAA28;
	input DATAA27;
	input DATAA26;
	input DATAA25;
	input DATAA24;
	input DATAA23;
	input DATAA22;
	input DATAA21;
	input DATAA20;
	input DATAA19;
	input DATAA18;
	input DATAA17;
	input DATAA16;
	input DATAA15;
	input DATAA14;
	input DATAA13;
	input DATAA12;
	input DATAA11;
	input DATAA10;
	input DATAA9;
	input DATAA8;
	input DATAA7;
	input DATAA6;
	input DATAA5;
	input DATAA4;
	input DATAA3;
	input DATAA2;
	input DATAA1;
	input DATAA0;
	input DATAB31;
	input DATAB30;
	input DATAB29;
	input DATAB28;
	input DATAB27;
	input DATAB26;
	input DATAB25;
	input DATAB24;
	input DATAB23;
	input DATAB22;
	input DATAB21;
	input DATAB20;
	input DATAB19;
	input DATAB18;
	input DATAB17;
	input DATAB16;
	input DATAB15;
	input DATAB14;
	input DATAB13;
	input DATAB12;
	input DATAB11;
	input DATAB10;
	input DATAB9;
	input DATAB8;
	input DATAB7;
	input DATAB6;
	input DATAB5;
	input DATAB4;
	input DATAB3;
	input DATAB2;
	input DATAB1;
	input DATAB0;
	input DATAC4;
	input DATAC3;
	input DATAC2;
	input DATAC1;
	input DATAC0;
	input OPC6;
	input OPC5;
	input OPC4;
	input OPC3;
	input OPC2;
	input OPC1;
	input OPC0;
	input OPCCUSTOM;
	input RADDRA4;
	input RADDRA3;
	input RADDRA2;
	input RADDRA1;
	input RADDRA0;
	input RADDRB4;
	input RADDRB3;
	input RADDRB2;
	input RADDRB1;
	input RADDRB0;
	output RDATAA31;
	output RDATAA30;
	output RDATAA29;
	output RDATAA28;
	output RDATAA27;
	output RDATAA26;
	output RDATAA25;
	output RDATAA24;
	output RDATAA23;
	output RDATAA22;
	output RDATAA21;
	output RDATAA20;
	output RDATAA19;
	output RDATAA18;
	output RDATAA17;
	output RDATAA16;
	output RDATAA15;
	output RDATAA14;
	output RDATAA13;
	output RDATAA12;
	output RDATAA11;
	output RDATAA10;
	output RDATAA9;
	output RDATAA8;
	output RDATAA7;
	output RDATAA6;
	output RDATAA5;
	output RDATAA4;
	output RDATAA3;
	output RDATAA2;
	output RDATAA1;
	output RDATAA0;
	output RDATAB31;
	output RDATAB30;
	output RDATAB29;
	output RDATAB28;
	output RDATAB27;
	output RDATAB26;
	output RDATAB25;
	output RDATAB24;
	output RDATAB23;
	output RDATAB22;
	output RDATAB21;
	output RDATAB20;
	output RDATAB19;
	output RDATAB18;
	output RDATAB17;
	output RDATAB16;
	output RDATAB15;
	output RDATAB14;
	output RDATAB13;
	output RDATAB12;
	output RDATAB11;
	output RDATAB10;
	output RDATAB9;
	output RDATAB8;
	output RDATAB7;
	output RDATAB6;
	output RDATAB5;
	output RDATAB4;
	output RDATAB3;
	output RDATAB2;
	output RDATAB1;
	output RDATAB0;
	input REGCLK;
	input REGCLKEN;
	input REGRST;
	output RESULT31;
	output RESULT30;
	output RESULT29;
	output RESULT28;
	output RESULT27;
	output RESULT26;
	output RESULT25;
	output RESULT24;
	output RESULT23;
	output RESULT22;
	output RESULT21;
	output RESULT20;
	output RESULT19;
	output RESULT18;
	output RESULT17;
	output RESULT16;
	output RESULT15;
	output RESULT14;
	output RESULT13;
	output RESULT12;
	output RESULT11;
	output RESULT10;
	output RESULT9;
	output RESULT8;
	output RESULT7;
	output RESULT6;
	output RESULT5;
	output RESULT4;
	output RESULT3;
	output RESULT2;
	output RESULT1;
	output RESULT0;
	input SCANCLK;
	input SCANRST;
	input WADDR4;
	input WADDR3;
	input WADDR2;
	input WADDR1;
	input WADDR0;
	input WDROTATE1;
	input WDROTATE0;
	input WDSIGNEXT;
	input WDSIZE1;
	input WDSIZE0;
	input WDATA31;
	input WDATA30;
	input WDATA29;
	input WDATA28;
	input WDATA27;
	input WDATA26;
	input WDATA25;
	input WDATA24;
	input WDATA23;
	input WDATA22;
	input WDATA21;
	input WDATA20;
	input WDATA19;
	input WDATA18;
	input WDATA17;
	input WDATA16;
	input WDATA15;
	input WDATA14;
	input WDATA13;
	input WDATA12;
	input WDATA11;
	input WDATA10;
	input WDATA9;
	input WDATA8;
	input WDATA7;
	input WDATA6;
	input WDATA5;
	input WDATA4;
	input WDATA3;
	input WDATA2;
	input WDATA1;
	input WDATA0;
	input WREN;

	parameter ALURST_ACTIVELOW = "DISABLE";
	parameter GSR = "ENABLED";
	parameter INREG = "DISABLE";
	parameter MULFXP_ROUND = "ENABLE";
	parameter OUTREG = "DISABLE";
	parameter REGRST_ACTIVELOW = "DISABLE";
	parameter RETAIN = "ENABLE";
	parameter RFASYNC_RD = "SYNC_RD";
	parameter RFR0_RO = "R0READONLY";
	parameter RFUNALIA_WR = "DISABLE";
	parameter RFWCLK_INV = "SIG";

endmodule

module BNKREF18_CORE (STDBYINR, STDBYDIF, PVTSNKI6, PVTSNKI5, PVTSNKI4, PVTSNKI3, PVTSNKI2, PVTSNKI1, PVTSNKI0, PVTSRCI6, PVTSRCI5, PVTSRCI4, PVTSRCI3, PVTSRCI2, PVTSRCI1, PVTSRCI0, PVTCODE6, PVTCODE5, PVTCODE4, PVTCODE3, PVTCODE2, PVTCODE1, PVTCODE0, PVTSEL); //synthesis syn_black_box syn_noprune=1 syn_lib_cell=1

	input STDBYINR;
	input STDBYDIF;
	input PVTSNKI6;
	input PVTSNKI5;
	input PVTSNKI4;
	input PVTSNKI3;
	input PVTSNKI2;
	input PVTSNKI1;
	input PVTSNKI0;
	input PVTSRCI6;
	input PVTSRCI5;
	input PVTSRCI4;
	input PVTSRCI3;
	input PVTSRCI2;
	input PVTSRCI1;
	input PVTSRCI0;
	output PVTCODE6;
	output PVTCODE5;
	output PVTCODE4;
	output PVTCODE3;
	output PVTCODE2;
	output PVTCODE1;
	output PVTCODE0;
	input PVTSEL;

	parameter BANK = "0b0000";
	parameter STANDBY_DIFFIO = "DISABLED";
	parameter STANDBY_INR = "DISABLED";

endmodule

module BNKREF33_CORE (PVTSEL, PVTSNKI6, PVTSNKI5, PVTSNKI4, PVTSNKI3, PVTSNKI2, PVTSNKI1, PVTSNKI0, PVTSRCI6, PVTSRCI5, PVTSRCI4, PVTSRCI3, PVTSRCI2, PVTSRCI1, PVTSRCI0, PVTCODE6, PVTCODE5, PVTCODE4, PVTCODE3, PVTCODE2, PVTCODE1, PVTCODE0); //synthesis syn_black_box syn_lib_cell=1

	input PVTSEL;
	input PVTSNKI6;
	input PVTSNKI5;
	input PVTSNKI4;
	input PVTSNKI3;
	input PVTSNKI2;
	input PVTSNKI1;
	input PVTSNKI0;
	input PVTSRCI6;
	input PVTSRCI5;
	input PVTSRCI4;
	input PVTSRCI3;
	input PVTSRCI2;
	input PVTSRCI1;
	input PVTSRCI0;
	output PVTCODE6;
	output PVTCODE5;
	output PVTCODE4;
	output PVTCODE3;
	output PVTCODE2;
	output PVTCODE1;
	output PVTCODE0;

	parameter BANK = "0b0000";

endmodule

module DIFFIO18_CORE (I, DOLP, B, O, INLP, T, INADC, HSRXEN, HSTXEN); //synthesis syn_black_box black_box_pad_pin="B" syn_lib_cell=1

	input I;
	input DOLP;
	inout B;
	output O;
	output INLP;
	input T;
	output INADC;
	input HSRXEN;
	input HSTXEN;

	parameter MIPI_ID = "0";
	parameter PULLMODE = "DOWN";
	parameter ENADC_IN = "DISABLED";
	parameter MIPI = "DISABLED";

endmodule

module CONFIG_CLKRST_CORE (HSE_CLK, JTAG_LRST_N, LMMI_CLK, LMMI_CLK_O, LMMI_LRST_N, LMMI_RST, MBISTCLK, OSCCLK, SEDC_CLK, SEDC_LRST_N, SEDC_RST, CFG_CLK, SMCLK_RST, WDT_CLK, WDT_LRST_N, WDT_RST); //synthesis syn_black_box syn_lib_cell=1

	output HSE_CLK;
	input JTAG_LRST_N;
	input LMMI_CLK;
	output LMMI_CLK_O;
	input LMMI_LRST_N;
	output LMMI_RST;
    input MBISTCLK;
	input OSCCLK;
	input SEDC_CLK;
	input SEDC_LRST_N;
	output SEDC_RST;
	output CFG_CLK;
	output SMCLK_RST;
	output WDT_CLK;
	input WDT_LRST_N;
	output WDT_RST;

	parameter MCJTAGGSRNDIS = "EN";
	parameter MCLMMIGSRNDIS = "EN";
	parameter MCSEDCGSRNDIS = "EN";
	parameter MCWDTGSRNDIS = "EN";
	parameter SMCLK_DIV = "3";

endmodule




module CONFIG_JTAG_CORE (JCE1, JCE2, JRSTN, JRTI1, JRTI2, JSHIFT, JTDI, JUPDATE, JTDO1, JTDO2, SMCLK, TCK, JTCK, TDI, TDO_OEN, TDO, TMS); //synthesis syn_black_box syn_lib_cell=1

	output JCE1;
	output JCE2;
	output JRSTN;
	output JRTI1;
	output JRTI2;
	output JSHIFT;
	output JTDI;
	output JUPDATE;
	input JTDO1;
	input JTDO2;
	input SMCLK;
	input TCK;
	output JTCK;
	input TDI;
	output TDO_OEN;
	output TDO;
	input TMS;

	parameter MCER1EXIST = "NEXIST";
	parameter MCER2EXIST = "NEXIST";

endmodule

module CONFIG_LMMI_CORE (LMMIOFFSET7, LMMIOFFSET6, LMMIOFFSET5, LMMIOFFSET4, LMMIOFFSET3, LMMIOFFSET2, LMMIOFFSET1, LMMIOFFSET0, LMMICLK, LMMIRDATA7, LMMIRDATA6, LMMIRDATA5, LMMIRDATA4, LMMIRDATA3, LMMIRDATA2, LMMIRDATA1, LMMIRDATA0, LMMIRDATAVALID, LMMIREADY, LMMIRESETN, LMMIREQUEST, LMMIWDATA7, LMMIWDATA6, LMMIWDATA5, LMMIWDATA4, LMMIWDATA3, LMMIWDATA2, LMMIWDATA1, LMMIWDATA0, LMMIWRRDN, RSTSMCLK, SMCLK); //synthesis syn_black_box syn_lib_cell=1

	input LMMIOFFSET7;
	input LMMIOFFSET6;
	input LMMIOFFSET5;
	input LMMIOFFSET4;
	input LMMIOFFSET3;
	input LMMIOFFSET2;
	input LMMIOFFSET1;
	input LMMIOFFSET0;
	input LMMICLK;
	output LMMIRDATA7;
	output LMMIRDATA6;
	output LMMIRDATA5;
	output LMMIRDATA4;
	output LMMIRDATA3;
	output LMMIRDATA2;
	output LMMIRDATA1;
	output LMMIRDATA0;
	output LMMIRDATAVALID;
	output LMMIREADY;
	input LMMIRESETN;
	input LMMIREQUEST;
	input LMMIWDATA7;
	input LMMIWDATA6;
	input LMMIWDATA5;
	input LMMIWDATA4;
	input LMMIWDATA3;
	input LMMIWDATA2;
	input LMMIWDATA1;
	input LMMIWDATA0;
	input LMMIWRRDN;
	input RSTSMCLK;
	input SMCLK;

	parameter LMMI_EN = "DIS";

endmodule

module CONFIG_MULTIBOOT_CORE (CIBAUTOREBOOT, CIBMSPIMADDR31, CIBMSPIMADDR30, CIBMSPIMADDR29, CIBMSPIMADDR28, CIBMSPIMADDR27, CIBMSPIMADDR26, CIBMSPIMADDR25, CIBMSPIMADDR24, CIBMSPIMADDR23, CIBMSPIMADDR22, CIBMSPIMADDR21, CIBMSPIMADDR20, CIBMSPIMADDR19, CIBMSPIMADDR18, CIBMSPIMADDR17, CIBMSPIMADDR16, CIBMSPIMADDR15, CIBMSPIMADDR14, CIBMSPIMADDR13, CIBMSPIMADDR12, CIBMSPIMADDR11, CIBMSPIMADDR10, CIBMSPIMADDR9, CIBMSPIMADDR8, CIBMSPIMADDR7, CIBMSPIMADDR6, CIBMSPIMADDR5, CIBMSPIMADDR4, CIBMSPIMADDR3, CIBMSPIMADDR2, CIBMSPIMADDR1, CIBMSPIMADDR0); //synthesis syn_black_box syn_noprune=1 syn_lib_cell=1

	input CIBAUTOREBOOT;
	input CIBMSPIMADDR31;
	input CIBMSPIMADDR30;
	input CIBMSPIMADDR29;
	input CIBMSPIMADDR28;
	input CIBMSPIMADDR27;
	input CIBMSPIMADDR26;
	input CIBMSPIMADDR25;
	input CIBMSPIMADDR24;
	input CIBMSPIMADDR23;
	input CIBMSPIMADDR22;
	input CIBMSPIMADDR21;
	input CIBMSPIMADDR20;
	input CIBMSPIMADDR19;
	input CIBMSPIMADDR18;
	input CIBMSPIMADDR17;
	input CIBMSPIMADDR16;
	input CIBMSPIMADDR15;
	input CIBMSPIMADDR14;
	input CIBMSPIMADDR13;
	input CIBMSPIMADDR12;
	input CIBMSPIMADDR11;
	input CIBMSPIMADDR10;
	input CIBMSPIMADDR9;
	input CIBMSPIMADDR8;
	input CIBMSPIMADDR7;
	input CIBMSPIMADDR6;
	input CIBMSPIMADDR5;
	input CIBMSPIMADDR4;
	input CIBMSPIMADDR3;
	input CIBMSPIMADDR2;
	input CIBMSPIMADDR1;
	input CIBMSPIMADDR0;

	parameter MSPIADDR = "0b00000000000000000000000000000000";
	parameter SOURCESEL = "DIS";

endmodule

module CONFIG_SEDC_CORE (CIBSED1ENABLE, CIBSEDCCOF, CIBSEDCENABLE, CIBSEDCMODE, CIBSEDCSTART, OSCCLKSEDC, RSTSEDC, SEDCBUSYCIB, SEDCDSRERRLOCCIB12, SEDCDSRERRLOCCIB11, SEDCDSRERRLOCCIB10, SEDCDSRERRLOCCIB9, SEDCDSRERRLOCCIB8, SEDCDSRERRLOCCIB7, SEDCDSRERRLOCCIB6, SEDCDSRERRLOCCIB5, SEDCDSRERRLOCCIB4, SEDCDSRERRLOCCIB3, SEDCDSRERRLOCCIB2, SEDCDSRERRLOCCIB1, SEDCDSRERRLOCCIB0, SEDCERR1CIB, SEDCERRCCIB, SEDCERRCRCCIB, SEDCERRMCIB, SEDCFRMERRLOCCIB15, SEDCFRMERRLOCCIB14, SEDCFRMERRLOCCIB13, SEDCFRMERRLOCCIB12, SEDCFRMERRLOCCIB11, SEDCFRMERRLOCCIB10, SEDCFRMERRLOCCIB9, SEDCFRMERRLOCCIB8, SEDCFRMERRLOCCIB7, SEDCFRMERRLOCCIB6, SEDCFRMERRLOCCIB5, SEDCFRMERRLOCCIB4, SEDCFRMERRLOCCIB3, SEDCFRMERRLOCCIB2, SEDCFRMERRLOCCIB1, SEDCFRMERRLOCCIB0); //synthesis syn_black_box syn_lib_cell=1

	input CIBSED1ENABLE;
	input CIBSEDCCOF;
	input CIBSEDCENABLE;
	input CIBSEDCMODE;
	input CIBSEDCSTART;
	input OSCCLKSEDC;
	input RSTSEDC;
	output SEDCBUSYCIB;
	output SEDCDSRERRLOCCIB12;
	output SEDCDSRERRLOCCIB11;
	output SEDCDSRERRLOCCIB10;
	output SEDCDSRERRLOCCIB9;
	output SEDCDSRERRLOCCIB8;
	output SEDCDSRERRLOCCIB7;
	output SEDCDSRERRLOCCIB6;
	output SEDCDSRERRLOCCIB5;
	output SEDCDSRERRLOCCIB4;
	output SEDCDSRERRLOCCIB3;
	output SEDCDSRERRLOCCIB2;
	output SEDCDSRERRLOCCIB1;
	output SEDCDSRERRLOCCIB0;
	output SEDCERR1CIB;
	output SEDCERRCCIB;
	output SEDCERRCRCCIB;
	output SEDCERRMCIB;
	output SEDCFRMERRLOCCIB15;
	output SEDCFRMERRLOCCIB14;
	output SEDCFRMERRLOCCIB13;
	output SEDCFRMERRLOCCIB12;
	output SEDCFRMERRLOCCIB11;
	output SEDCFRMERRLOCCIB10;
	output SEDCFRMERRLOCCIB9;
	output SEDCFRMERRLOCCIB8;
	output SEDCFRMERRLOCCIB7;
	output SEDCFRMERRLOCCIB6;
	output SEDCFRMERRLOCCIB5;
	output SEDCFRMERRLOCCIB4;
	output SEDCFRMERRLOCCIB3;
	output SEDCFRMERRLOCCIB2;
	output SEDCFRMERRLOCCIB1;
	output SEDCFRMERRLOCCIB0;

	parameter SEDCEN = "DIS";

endmodule

module CONFIG_WDT_CORE (CIBWDTRELOAD, WDT_CLK, WDT_RST); //synthesis syn_black_box syn_noprune=1 syn_lib_cell=1

	input CIBWDTRELOAD;
	input WDT_CLK;
	input WDT_RST;

	parameter WDTEN = "DIS";
	parameter WDTMODE = "SINGLE";
	parameter WDTVALUE = "0b000000000000000000";

endmodule

module DDRDLL_CORE (CODE8, CODE7, CODE6, CODE5, CODE4, CODE3, CODE2, CODE1, CODE0, FREEZE, LOCK, CLKIN, RST, DCNTL8, DCNTL7, DCNTL6, DCNTL5, DCNTL4, DCNTL3, DCNTL2, DCNTL1, DCNTL0, UDDCNTL_N); //synthesis syn_black_box syn_lib_cell=1

	output CODE8;
	output CODE7;
	output CODE6;
	output CODE5;
	output CODE4;
	output CODE3;
	output CODE2;
	output CODE1;
	output CODE0;
	input FREEZE;
	output LOCK;
	input CLKIN;
	input RST;
	output DCNTL8;
	output DCNTL7;
	output DCNTL6;
	output DCNTL5;
	output DCNTL4;
	output DCNTL3;
	output DCNTL2;
	output DCNTL1;
	output DCNTL0;
	input UDDCNTL_N;

	parameter GSR = "ENABLED";
	parameter ENA_ROUNDOFF = "ENABLED";
	parameter FORCE_MAX_DELAY = "CODE_OR_LOCK_FROM_DLL_LOOP";

endmodule

module DLLDEL_CORE (CLKIN, CLKOUT, CODE8, CODE7, CODE6, CODE5, CODE4, CODE3, CODE2, CODE1, CODE0, COUT, DIR, LOAD_N, MOVE); //synthesis syn_black_box syn_lib_cell=1

	input CLKIN;
	output CLKOUT;
	input CODE8;
	input CODE7;
	input CODE6;
	input CODE5;
	input CODE4;
	input CODE3;
	input CODE2;
	input CODE1;
	input CODE0;
	output COUT;
	input DIR;
	input LOAD_N;
	input MOVE;

	parameter ADJUST = "0";
	parameter DEL_ADJUST = "PLUS";
	parameter ENABLE = "DISABLED";

endmodule

module DPHY_CORE (BITCKEXT, CKN, CKP, CLKREF, D0ACTIVE1, D0ACTIVE0, D0BYTCNT9, D0BYTCNT8, D0BYTCNT7, D0BYTCNT6, D0BYTCNT5, D0BYTCNT4, D0BYTCNT3, D0BYTCNT2, D0BYTCNT1, D0BYTCNT0, D0ERRCNT9, D0ERRCNT8, D0ERRCNT7, D0ERRCNT6, D0ERRCNT5, D0ERRCNT4, D0ERRCNT3, D0ERRCNT2, D0ERRCNT1, D0ERRCNT0, D0PASS1, D0PASS0, D0VALID1, D0VALID0, D1ACTIVE1, D1ACTIVE0, D1BYTCNT9, D1BYTCNT8, D1BYTCNT7, D1BYTCNT6, D1BYTCNT5, D1BYTCNT4, D1BYTCNT3, D1BYTCNT2, D1BYTCNT1, D1BYTCNT0, D1ERRCNT9, D1ERRCNT8, D1ERRCNT7, D1ERRCNT6, D1ERRCNT5, D1ERRCNT4, D1ERRCNT3, D1ERRCNT2, D1ERRCNT1, D1ERRCNT0, D1PASS1, D1PASS0, D1VALID1, D1VALID0, D2ACTIVE1, D2ACTIVE0, D2BYTCNT9, D2BYTCNT8, D2BYTCNT7, D2BYTCNT6, D2BYTCNT5, D2BYTCNT4, D2BYTCNT3, D2BYTCNT2, D2BYTCNT1, D2BYTCNT0, D2ERRCNT9, D2ERRCNT8, D2ERRCNT7, D2ERRCNT6, D2ERRCNT5, D2ERRCNT4, D2ERRCNT3, D2ERRCNT2, D2ERRCNT1, D2ERRCNT0, D2PASS1, D2PASS0, D2VALID1, D2VALID0, D3ACTIVE1, D3ACTIVE0, D3BYTCNT9, D3BYTCNT8, D3BYTCNT7, D3BYTCNT6, D3BYTCNT5, D3BYTCNT4, D3BYTCNT3, D3BYTCNT2, D3BYTCNT1, D3BYTCNT0, D3ERRCNT9, D3ERRCNT8, D3ERRCNT7, D3ERRCNT6, D3ERRCNT5, D3ERRCNT4, D3ERRCNT3, D3ERRCNT2, D3ERRCNT1, D3ERRCNT0, D3PASS1, D3PASS0, D3VALID1, D3VALID0, DCTSTOUT9, DCTSTOUT8, DCTSTOUT7, DCTSTOUT6, DCTSTOUT5, DCTSTOUT4, DCTSTOUT3, DCTSTOUT2, DCTSTOUT1, DCTSTOUT0, DN0, DN1, DN2, DN3, DP0, DP1, DP2, DP3, LOCK, PDDPHY, PDPLL, SCCLKIN, SCRSTNIN, UDIR, UED0THEN, UERCLP0, UERCLP1, UERCTRL, UERE, UERSTHS, UERSSHS, UERSE, UFRXMODE, UTXMDTX, URXACTHS, URXCKE, URXCKINE, URXDE7, URXDE6, URXDE5, URXDE4, URXDE3, URXDE2, URXDE1, URXDE0, URXDHS15, URXDHS14, URXDHS13, URXDHS12, URXDHS11, URXDHS10, URXDHS9, URXDHS8, URXDHS7, URXDHS6, URXDHS5, URXDHS4, URXDHS3, URXDHS2, URXDHS1, URXDHS0, URXLPDTE, URXSKCHS, URXDRX, URXSHS3, URXSHS2, URXSHS1, URXSHS0, URE0D3DP, URE1D3DN, URE2CKDP, URE3CKDN, URXULPSE, URXVDE, URXVDHS3, URXVDHS2, URXVDHS1, URXVDHS0, USSTT, UTDIS, UTXCKE, UDE0D0TN, UDE1D1TN, UDE2D2TN, UDE3D3TN, UDE4CKTN, UDE5D0RN, UDE6D1RN, UDE7D2RN, UTXDHS31, UTXDHS30, UTXDHS29, UTXDHS28, UTXDHS27, UTXDHS26, UTXDHS25, UTXDHS24, UTXDHS23, UTXDHS22, UTXDHS21, UTXDHS20, UTXDHS19, UTXDHS18, UTXDHS17, UTXDHS16, UTXDHS15, UTXDHS14, UTXDHS13, UTXDHS12, UTXDHS11, UTXDHS10, UTXDHS9, UTXDHS8, UTXDHS7, UTXDHS6, UTXDHS5, UTXDHS4, UTXDHS3, UTXDHS2, UTXDHS1, UTXDHS0, UTXENER, UTXRRS, UTXRYP, UTXRYSK, UTXRD0EN, UTRD0SEN, UTXSKD0N, UTXTGE0, UTXTGE1, UTXTGE2, UTXTGE3, UTXULPSE, UTXUPSEX, UTXVDE, UTXWVDHS3, UTXWVDHS2, UTXWVDHS1, UTXWVDHS0, UUSAN, U1DIR, U1ENTHEN, U1ERCLP0, U1ERCLP1, U1ERCTRL, U1ERE, U1ERSTHS, U1ERSSHS, U1ERSE, U1FRXMD, U1FTXST, U1RXATHS, U1RXCKE, U1RXDE7, U1RXDE6, U1RXDE5, U1RXDE4, U1RXDE3, U1RXDE2, U1RXDE1, U1RXDE0, U1RXDHS15, U1RXDHS14, U1RXDHS13, U1RXDHS12, U1RXDHS11, U1RXDHS10, U1RXDHS9, U1RXDHS8, U1RXDHS7, U1RXDHS6, U1RXDHS5, U1RXDHS4, U1RXDHS3, U1RXDHS2, U1RXDHS1, U1RXDHS0, U1RXDTE, U1RXSKS, U1RXSK, U1RXSHS3, U1RXSHS2, U1RXSHS1, U1RXSHS0, U1RE0D, U1RE1CN, U1RE2D, U1RE3N, U1RXUPSE, U1RXVDE, U1RXVDHS3, U1RXVDHS2, U1RXVDHS1, U1RXVDHS0, U1SSTT, U1TDIS, U1TREQ, U1TDE0D3, U1TDE1CK, U1TDE2D0, U1TDE3D1, U1TDE4D2, U1TDE5D3, U1TDE6, U1TDE7, U1TXDHS31, U1TXDHS30, U1TXDHS29, U1TXDHS28, U1TXDHS27, U1TXDHS26, U1TXDHS25, U1TXDHS24, U1TXDHS23, U1TXDHS22, U1TXDHS21, U1TXDHS20, U1TXDHS19, U1TXDHS18, U1TXDHS17, U1TXDHS16, U1TXDHS15, U1TXDHS14, U1TXDHS13, U1TXDHS12, U1TXDHS11, U1TXDHS10, U1TXDHS9, U1TXDHS8, U1TXDHS7, U1TXDHS6, U1TXDHS5, U1TXDHS4, U1TXDHS3, U1TXDHS2, U1TXDHS1, U1TXDHS0, U1TXLPD, U1TXRYE, U1TXRY, U1TXRYSK, U1TXREQ, U1TXREQH, U1TXSK, U1TXTGE0, U1TXTGE1, U1TXTGE2, U1TXTGE3, U1TXUPSE, U1TXUPSX, U1TXVDE, U1TXWVHS3, U1TXWVHS2, U1TXWVHS1, U1TXWVHS0, U1USAN, U2DIR, U2END2, U2ERCLP0, U2ERCLP1, U2ERCTRL, U2ERE, U2ERSTHS, U2ERSSHS, U2ERSE, U2FRXMD, U2FTXST, U2RXACHS, U2RXCKE, U2RXDE7, U2RXDE6, U2RXDE5, U2RXDE4, U2RXDE3, U2RXDE2, U2RXDE1, U2RXDE0, U2RXDHS15, U2RXDHS14, U2RXDHS13, U2RXDHS12, U2RXDHS11, U2RXDHS10, U2RXDHS9, U2RXDHS8, U2RXDHS7, U2RXDHS6, U2RXDHS5, U2RXDHS4, U2RXDHS3, U2RXDHS2, U2RXDHS1, U2RXDHS0, U2RPDTE, U2RXSK, U2RXSKC, U2RXSHS3, U2RXSHS2, U2RXSHS1, U2RXSHS0, U2RE0D2, U2RE1D2, U2RE2D3, U2RE3D3, U2RXUPSE, U2RXVDE, U2RXVDHS3, U2RXVDHS2, U2RXVDHS1, U2RXVDHS0, U2SSTT, U2TDIS, U2TREQ, U2TDE0D0, U2TDE1D1, U2TDE2D2, U2TDE3D3, U2TDE4CK, U2TDE5D0, U2TDE6D1, U2TDE7D2, U2TXDHS31, U2TXDHS30, U2TXDHS29, U2TXDHS28, U2TXDHS27, U2TXDHS26, U2TXDHS25, U2TXDHS24, U2TXDHS23, U2TXDHS22, U2TXDHS21, U2TXDHS20, U2TXDHS19, U2TXDHS18, U2TXDHS17, U2TXDHS16, U2TXDHS15, U2TXDHS14, U2TXDHS13, U2TXDHS12, U2TXDHS11, U2TXDHS10, U2TXDHS9, U2TXDHS8, U2TXDHS7, U2TXDHS6, U2TXDHS5, U2TXDHS4, U2TXDHS3, U2TXDHS2, U2TXDHS1, U2TXDHS0, U2TPDTE, U2TXRYE, U2TXRYH, U2TXRYSK, U2TXREQ, U2TXREQH, U2TXSKC, U2TXTGE0, U2TXTGE1, U2TXTGE2, U2TXTGE3, U2TXUPSE, U2TXUPSX, U2TXVDE, U2TXWVHS3, U2TXWVHS2, U2TXWVHS1, U2TXWVHS0, U2USAN, U3DIR, U3END3, U3ERCLP0, U3ERCLP1, U3ERCTRL, U3ERE, U3ERSTHS, U3ERSSHS, U3ERSE, U3FRXMD, U3FTXST, U3RXATHS, U3RXCKE, U3RXDE7, U3RXDE6, U3RXDE5, U3RXDE4, U3RXDE3, U3RXDE2, U3RXDE1, U3RXDE0, U3RXDHS15, U3RXDHS14, U3RXDHS13, U3RXDHS12, U3RXDHS11, U3RXDHS10, U3RXDHS9, U3RXDHS8, U3RXDHS7, U3RXDHS6, U3RXDHS5, U3RXDHS4, U3RXDHS3, U3RXDHS2, U3RXDHS1, U3RXDHS0, U3RPDTE, U3RXSK, U3RXSKC, U3RXSHS3, U3RXSHS2, U3RXSHS1, U3RXSHS0, U3RE0CK, U3RE1CK, U3RE2, U3RE3, U3RXUPSE, U3RXVDE, U3RXVDHS3, U3RXVDHS2, U3RXVDHS1, U3RXVDHS0, U3SSTT, U3TDISD2, U3TREQD2, U3TDE0D3, U3TDE1D0, U3TDE2D1, U3TDE3D2, U3TDE4D3, U3TDE5CK, U3TDE6, U3TDE7, U3TXDHS31, U3TXDHS30, U3TXDHS29, U3TXDHS28, U3TXDHS27, U3TXDHS26, U3TXDHS25, U3TXDHS24, U3TXDHS23, U3TXDHS22, U3TXDHS21, U3TXDHS20, U3TXDHS19, U3TXDHS18, U3TXDHS17, U3TXDHS16, U3TXDHS15, U3TXDHS14, U3TXDHS13, U3TXDHS12, U3TXDHS11, U3TXDHS10, U3TXDHS9, U3TXDHS8, U3TXDHS7, U3TXDHS6, U3TXDHS5, U3TXDHS4, U3TXDHS3, U3TXDHS2, U3TXDHS1, U3TXDHS0, U3TXLPDT, U3TXRY, U3TXRYHS, U3TXRYSK, U3TXREQ, U3TXREQH, U3TXSKC, U3TXTGE0, U3TXTGE1, U3TXTGE2, U3TXTGE3, U3TXULPS, U3TXUPSX, U3TXVD3, U3TXWVHS3, U3TXWVHS2, U3TXWVHS1, U3TXWVHS0, U3USAN, UCENCK, UCRXCKAT, UCRXUCKN, UCSSTT, UCTXREQH, UCTXUPSC, UCTXUPSX, UCUSAN, SCANCLK, SCANRST, LMMICLK, LMMIOFFSET4, LMMIOFFSET3, LMMIOFFSET2, LMMIOFFSET1, LMMIOFFSET0, LMMIRDATA3, LMMIRDATA2, LMMIRDATA1, LMMIRDATA0, LMMIRDATAVALID, LMMIREADY, LMMIREQUEST, LMMIRESETN, LMMIWDATA3, LMMIWDATA2, LMMIWDATA1, LMMIWDATA0, LMMIWRRDN, LTSTEN, LTSTLANE1, LTSTLANE0, URWDCKHS, UTRNREQ, UTWDCKHS, UCRXWCHS, OPCGLDCK, CLKLBACT); //synthesis syn_black_box black_box_pad_pin="CKN,CKP,DN0,DN1,DN2,DN3,DP0,DP1,DP2,DP3" syn_lib_cell=1

	input BITCKEXT;
	inout CKN;
	inout CKP;
	input CLKREF;
	output D0ACTIVE1;
	output D0ACTIVE0;
	output D0BYTCNT9;
	output D0BYTCNT8;
	output D0BYTCNT7;
	output D0BYTCNT6;
	output D0BYTCNT5;
	output D0BYTCNT4;
	output D0BYTCNT3;
	output D0BYTCNT2;
	output D0BYTCNT1;
	output D0BYTCNT0;
	output D0ERRCNT9;
	output D0ERRCNT8;
	output D0ERRCNT7;
	output D0ERRCNT6;
	output D0ERRCNT5;
	output D0ERRCNT4;
	output D0ERRCNT3;
	output D0ERRCNT2;
	output D0ERRCNT1;
	output D0ERRCNT0;
	output D0PASS1;
	output D0PASS0;
	output D0VALID1;
	output D0VALID0;
	output D1ACTIVE1;
	output D1ACTIVE0;
	output D1BYTCNT9;
	output D1BYTCNT8;
	output D1BYTCNT7;
	output D1BYTCNT6;
	output D1BYTCNT5;
	output D1BYTCNT4;
	output D1BYTCNT3;
	output D1BYTCNT2;
	output D1BYTCNT1;
	output D1BYTCNT0;
	output D1ERRCNT9;
	output D1ERRCNT8;
	output D1ERRCNT7;
	output D1ERRCNT6;
	output D1ERRCNT5;
	output D1ERRCNT4;
	output D1ERRCNT3;
	output D1ERRCNT2;
	output D1ERRCNT1;
	output D1ERRCNT0;
	output D1PASS1;
	output D1PASS0;
	output D1VALID1;
	output D1VALID0;
	output D2ACTIVE1;
	output D2ACTIVE0;
	output D2BYTCNT9;
	output D2BYTCNT8;
	output D2BYTCNT7;
	output D2BYTCNT6;
	output D2BYTCNT5;
	output D2BYTCNT4;
	output D2BYTCNT3;
	output D2BYTCNT2;
	output D2BYTCNT1;
	output D2BYTCNT0;
	output D2ERRCNT9;
	output D2ERRCNT8;
	output D2ERRCNT7;
	output D2ERRCNT6;
	output D2ERRCNT5;
	output D2ERRCNT4;
	output D2ERRCNT3;
	output D2ERRCNT2;
	output D2ERRCNT1;
	output D2ERRCNT0;
	output D2PASS1;
	output D2PASS0;
	output D2VALID1;
	output D2VALID0;
	output D3ACTIVE1;
	output D3ACTIVE0;
	output D3BYTCNT9;
	output D3BYTCNT8;
	output D3BYTCNT7;
	output D3BYTCNT6;
	output D3BYTCNT5;
	output D3BYTCNT4;
	output D3BYTCNT3;
	output D3BYTCNT2;
	output D3BYTCNT1;
	output D3BYTCNT0;
	output D3ERRCNT9;
	output D3ERRCNT8;
	output D3ERRCNT7;
	output D3ERRCNT6;
	output D3ERRCNT5;
	output D3ERRCNT4;
	output D3ERRCNT3;
	output D3ERRCNT2;
	output D3ERRCNT1;
	output D3ERRCNT0;
	output D3PASS1;
	output D3PASS0;
	output D3VALID1;
	output D3VALID0;
	output DCTSTOUT9;
	output DCTSTOUT8;
	output DCTSTOUT7;
	output DCTSTOUT6;
	output DCTSTOUT5;
	output DCTSTOUT4;
	output DCTSTOUT3;
	output DCTSTOUT2;
	output DCTSTOUT1;
	output DCTSTOUT0;
	inout DN0;
	inout DN1;
	inout DN2;
	inout DN3;
	inout DP0;
	inout DP1;
	inout DP2;
	inout DP3;
	output LOCK;
	input PDDPHY;
	input PDPLL;
	input SCCLKIN;
	input SCRSTNIN;
	output UDIR;
	input UED0THEN;
	output UERCLP0;
	output UERCLP1;
	output UERCTRL;
	output UERE;
	output UERSTHS;
	output UERSSHS;
	output UERSE;
	input UFRXMODE;
	input UTXMDTX;
	output URXACTHS;
	output URXCKE;
	input URXCKINE;
	output URXDE7;
	output URXDE6;
	output URXDE5;
	output URXDE4;
	output URXDE3;
	output URXDE2;
	output URXDE1;
	output URXDE0;
	output URXDHS15;
	output URXDHS14;
	output URXDHS13;
	output URXDHS12;
	output URXDHS11;
	output URXDHS10;
	output URXDHS9;
	output URXDHS8;
	output URXDHS7;
	output URXDHS6;
	output URXDHS5;
	output URXDHS4;
	output URXDHS3;
	output URXDHS2;
	output URXDHS1;
	output URXDHS0;
	output URXLPDTE;
	output URXSKCHS;
	output URXDRX;
	output URXSHS3;
	output URXSHS2;
	output URXSHS1;
	output URXSHS0;
	output URE0D3DP;
	output URE1D3DN;
	output URE2CKDP;
	output URE3CKDN;
	output URXULPSE;
	output URXVDE;
	output URXVDHS3;
	output URXVDHS2;
	output URXVDHS1;
	output URXVDHS0;
	output USSTT;
	input UTDIS;
	input UTXCKE;
	input UDE0D0TN;
	input UDE1D1TN;
	input UDE2D2TN;
	input UDE3D3TN;
	input UDE4CKTN;
	input UDE5D0RN;
	input UDE6D1RN;
	input UDE7D2RN;
	input UTXDHS31;
	input UTXDHS30;
	input UTXDHS29;
	input UTXDHS28;
	input UTXDHS27;
	input UTXDHS26;
	input UTXDHS25;
	input UTXDHS24;
	input UTXDHS23;
	input UTXDHS22;
	input UTXDHS21;
	input UTXDHS20;
	input UTXDHS19;
	input UTXDHS18;
	input UTXDHS17;
	input UTXDHS16;
	input UTXDHS15;
	input UTXDHS14;
	input UTXDHS13;
	input UTXDHS12;
	input UTXDHS11;
	input UTXDHS10;
	input UTXDHS9;
	input UTXDHS8;
	input UTXDHS7;
	input UTXDHS6;
	input UTXDHS5;
	input UTXDHS4;
	input UTXDHS3;
	input UTXDHS2;
	input UTXDHS1;
	input UTXDHS0;
	input UTXENER;
	output UTXRRS;
	output UTXRYP;
	output UTXRYSK;
	input UTXRD0EN;
	input UTRD0SEN;
	input UTXSKD0N;
	input UTXTGE0;
	input UTXTGE1;
	input UTXTGE2;
	input UTXTGE3;
	input UTXULPSE;
	input UTXUPSEX;
	input UTXVDE;
	input UTXWVDHS3;
	input UTXWVDHS2;
	input UTXWVDHS1;
	input UTXWVDHS0;
	output UUSAN;
	output U1DIR;
	input U1ENTHEN;
	output U1ERCLP0;
	output U1ERCLP1;
	output U1ERCTRL;
	output U1ERE;
	output U1ERSTHS;
	output U1ERSSHS;
	output U1ERSE;
	input U1FRXMD;
	input U1FTXST;
	output U1RXATHS;
	output U1RXCKE;
	output U1RXDE7;
	output U1RXDE6;
	output U1RXDE5;
	output U1RXDE4;
	output U1RXDE3;
	output U1RXDE2;
	output U1RXDE1;
	output U1RXDE0;
	output U1RXDHS15;
	output U1RXDHS14;
	output U1RXDHS13;
	output U1RXDHS12;
	output U1RXDHS11;
	output U1RXDHS10;
	output U1RXDHS9;
	output U1RXDHS8;
	output U1RXDHS7;
	output U1RXDHS6;
	output U1RXDHS5;
	output U1RXDHS4;
	output U1RXDHS3;
	output U1RXDHS2;
	output U1RXDHS1;
	output U1RXDHS0;
	output U1RXDTE;
	output U1RXSKS;
	output U1RXSK;
	output U1RXSHS3;
	output U1RXSHS2;
	output U1RXSHS1;
	output U1RXSHS0;
	output U1RE0D;
	output U1RE1CN;
	output U1RE2D;
	output U1RE3N;
	output U1RXUPSE;
	output U1RXVDE;
	output U1RXVDHS3;
	output U1RXVDHS2;
	output U1RXVDHS1;
	output U1RXVDHS0;
	output U1SSTT;
	input U1TDIS;
	input U1TREQ;
	input U1TDE0D3;
	input U1TDE1CK;
	input U1TDE2D0;
	input U1TDE3D1;
	input U1TDE4D2;
	input U1TDE5D3;
	input U1TDE6;
	input U1TDE7;
	input U1TXDHS31;
	input U1TXDHS30;
	input U1TXDHS29;
	input U1TXDHS28;
	input U1TXDHS27;
	input U1TXDHS26;
	input U1TXDHS25;
	input U1TXDHS24;
	input U1TXDHS23;
	input U1TXDHS22;
	input U1TXDHS21;
	input U1TXDHS20;
	input U1TXDHS19;
	input U1TXDHS18;
	input U1TXDHS17;
	input U1TXDHS16;
	input U1TXDHS15;
	input U1TXDHS14;
	input U1TXDHS13;
	input U1TXDHS12;
	input U1TXDHS11;
	input U1TXDHS10;
	input U1TXDHS9;
	input U1TXDHS8;
	input U1TXDHS7;
	input U1TXDHS6;
	input U1TXDHS5;
	input U1TXDHS4;
	input U1TXDHS3;
	input U1TXDHS2;
	input U1TXDHS1;
	input U1TXDHS0;
	input U1TXLPD;
	output U1TXRYE;
	output U1TXRY;
	output U1TXRYSK;
	input U1TXREQ;
	input U1TXREQH;
	input U1TXSK;
	input U1TXTGE0;
	input U1TXTGE1;
	input U1TXTGE2;
	input U1TXTGE3;
	input U1TXUPSE;
	input U1TXUPSX;
	input U1TXVDE;
	input U1TXWVHS3;
	input U1TXWVHS2;
	input U1TXWVHS1;
	input U1TXWVHS0;
	output U1USAN;
	output U2DIR;
	input U2END2;
	output U2ERCLP0;
	output U2ERCLP1;
	output U2ERCTRL;
	output U2ERE;
	output U2ERSTHS;
	output U2ERSSHS;
	output U2ERSE;
	input U2FRXMD;
	input U2FTXST;
	output U2RXACHS;
	output U2RXCKE;
	output U2RXDE7;
	output U2RXDE6;
	output U2RXDE5;
	output U2RXDE4;
	output U2RXDE3;
	output U2RXDE2;
	output U2RXDE1;
	output U2RXDE0;
	output U2RXDHS15;
	output U2RXDHS14;
	output U2RXDHS13;
	output U2RXDHS12;
	output U2RXDHS11;
	output U2RXDHS10;
	output U2RXDHS9;
	output U2RXDHS8;
	output U2RXDHS7;
	output U2RXDHS6;
	output U2RXDHS5;
	output U2RXDHS4;
	output U2RXDHS3;
	output U2RXDHS2;
	output U2RXDHS1;
	output U2RXDHS0;
	output U2RPDTE;
	output U2RXSK;
	output U2RXSKC;
	output U2RXSHS3;
	output U2RXSHS2;
	output U2RXSHS1;
	output U2RXSHS0;
	output U2RE0D2;
	output U2RE1D2;
	output U2RE2D3;
	output U2RE3D3;
	output U2RXUPSE;
	output U2RXVDE;
	output U2RXVDHS3;
	output U2RXVDHS2;
	output U2RXVDHS1;
	output U2RXVDHS0;
	output U2SSTT;
	input U2TDIS;
	input U2TREQ;
	input U2TDE0D0;
	input U2TDE1D1;
	input U2TDE2D2;
	input U2TDE3D3;
	input U2TDE4CK;
	input U2TDE5D0;
	input U2TDE6D1;
	input U2TDE7D2;
	input U2TXDHS31;
	input U2TXDHS30;
	input U2TXDHS29;
	input U2TXDHS28;
	input U2TXDHS27;
	input U2TXDHS26;
	input U2TXDHS25;
	input U2TXDHS24;
	input U2TXDHS23;
	input U2TXDHS22;
	input U2TXDHS21;
	input U2TXDHS20;
	input U2TXDHS19;
	input U2TXDHS18;
	input U2TXDHS17;
	input U2TXDHS16;
	input U2TXDHS15;
	input U2TXDHS14;
	input U2TXDHS13;
	input U2TXDHS12;
	input U2TXDHS11;
	input U2TXDHS10;
	input U2TXDHS9;
	input U2TXDHS8;
	input U2TXDHS7;
	input U2TXDHS6;
	input U2TXDHS5;
	input U2TXDHS4;
	input U2TXDHS3;
	input U2TXDHS2;
	input U2TXDHS1;
	input U2TXDHS0;
	input U2TPDTE;
	output U2TXRYE;
	output U2TXRYH;
	output U2TXRYSK;
	input U2TXREQ;
	input U2TXREQH;
	input U2TXSKC;
	input U2TXTGE0;
	input U2TXTGE1;
	input U2TXTGE2;
	input U2TXTGE3;
	input U2TXUPSE;
	input U2TXUPSX;
	input U2TXVDE;
	input U2TXWVHS3;
	input U2TXWVHS2;
	input U2TXWVHS1;
	input U2TXWVHS0;
	output U2USAN;
	output U3DIR;
	input U3END3;
	output U3ERCLP0;
	output U3ERCLP1;
	output U3ERCTRL;
	output U3ERE;
	output U3ERSTHS;
	output U3ERSSHS;
	output U3ERSE;
	input U3FRXMD;
	input U3FTXST;
	output U3RXATHS;
	output U3RXCKE;
	output U3RXDE7;
	output U3RXDE6;
	output U3RXDE5;
	output U3RXDE4;
	output U3RXDE3;
	output U3RXDE2;
	output U3RXDE1;
	output U3RXDE0;
	output U3RXDHS15;
	output U3RXDHS14;
	output U3RXDHS13;
	output U3RXDHS12;
	output U3RXDHS11;
	output U3RXDHS10;
	output U3RXDHS9;
	output U3RXDHS8;
	output U3RXDHS7;
	output U3RXDHS6;
	output U3RXDHS5;
	output U3RXDHS4;
	output U3RXDHS3;
	output U3RXDHS2;
	output U3RXDHS1;
	output U3RXDHS0;
	output U3RPDTE;
	output U3RXSK;
	output U3RXSKC;
	output U3RXSHS3;
	output U3RXSHS2;
	output U3RXSHS1;
	output U3RXSHS0;
	output U3RE0CK;
	output U3RE1CK;
	output U3RE2;
	output U3RE3;
	output U3RXUPSE;
	output U3RXVDE;
	output U3RXVDHS3;
	output U3RXVDHS2;
	output U3RXVDHS1;
	output U3RXVDHS0;
	output U3SSTT;
	input U3TDISD2;
	input U3TREQD2;
	input U3TDE0D3;
	input U3TDE1D0;
	input U3TDE2D1;
	input U3TDE3D2;
	input U3TDE4D3;
	input U3TDE5CK;
	input U3TDE6;
	input U3TDE7;
	input U3TXDHS31;
	input U3TXDHS30;
	input U3TXDHS29;
	input U3TXDHS28;
	input U3TXDHS27;
	input U3TXDHS26;
	input U3TXDHS25;
	input U3TXDHS24;
	input U3TXDHS23;
	input U3TXDHS22;
	input U3TXDHS21;
	input U3TXDHS20;
	input U3TXDHS19;
	input U3TXDHS18;
	input U3TXDHS17;
	input U3TXDHS16;
	input U3TXDHS15;
	input U3TXDHS14;
	input U3TXDHS13;
	input U3TXDHS12;
	input U3TXDHS11;
	input U3TXDHS10;
	input U3TXDHS9;
	input U3TXDHS8;
	input U3TXDHS7;
	input U3TXDHS6;
	input U3TXDHS5;
	input U3TXDHS4;
	input U3TXDHS3;
	input U3TXDHS2;
	input U3TXDHS1;
	input U3TXDHS0;
	input U3TXLPDT;
	output U3TXRY;
	output U3TXRYHS;
	output U3TXRYSK;
	input U3TXREQ;
	input U3TXREQH;
	input U3TXSKC;
	input U3TXTGE0;
	input U3TXTGE1;
	input U3TXTGE2;
	input U3TXTGE3;
	input U3TXULPS;
	input U3TXUPSX;
	input U3TXVD3;
	input U3TXWVHS3;
	input U3TXWVHS2;
	input U3TXWVHS1;
	input U3TXWVHS0;
	output U3USAN;
	input UCENCK;
	output UCRXCKAT;
	output UCRXUCKN;
	output UCSSTT;
	input UCTXREQH;
	input UCTXUPSC;
	input UCTXUPSX;
	output UCUSAN;
	input SCANCLK;
	input SCANRST;
	input LMMICLK;
	input LMMIOFFSET4;
	input LMMIOFFSET3;
	input LMMIOFFSET2;
	input LMMIOFFSET1;
	input LMMIOFFSET0;
	output LMMIRDATA3;
	output LMMIRDATA2;
	output LMMIRDATA1;
	output LMMIRDATA0;
	output LMMIRDATAVALID;
	output LMMIREADY;
	input LMMIREQUEST;
	input LMMIRESETN;
	input LMMIWDATA3;
	input LMMIWDATA2;
	input LMMIWDATA1;
	input LMMIWDATA0;
	input LMMIWRRDN;
	input LTSTEN;
	input LTSTLANE1;
	input LTSTLANE0;
	output URWDCKHS;
	input UTRNREQ;
	output UTWDCKHS;
	output UCRXWCHS;
	input OPCGLDCK;
	output CLKLBACT;

	parameter GSR = "ENABLED";
	parameter AUTO_PD_EN = "POWERED_UP";
	parameter CFG_NUM_LANES = "ONE_LANE";
	parameter CM = "0b00000000";
	parameter CN = "0b00000";
	parameter CO = "0b000";
	parameter CONT_CLK_MODE = "DISABLED";
	parameter DESKEW_EN = "DISABLED";
	parameter DSI_CSI = "CSI2_APP";
	parameter EN_CIL = "CIL_ENABLED";
	parameter HSEL = "DISABLED";
	parameter LANE0_SEL = "LANE_0";
	parameter LOCK_BYP = "GATE_TXBYTECLKHS";
	parameter MASTER_SLAVE = "SLAVE";
	parameter PLLCLKBYPASS = "REGISTERED";
	parameter RSEL = "0b00";
	parameter RXCDRP = "0b00";
	parameter RXDATAWIDTHHS = "0b00";
	parameter RXLPRP = "0b000";
	parameter TEST_ENBL = "0b000000";
	parameter TEST_PATTERN = "0b00000000000000000000000000000000";
	parameter TST = "0b1001";
	parameter TXDATAWIDTHHS = "0b00";
	parameter U_PRG_HS_PREPARE = "0b00";
	parameter U_PRG_HS_TRAIL = "0b000000";
	parameter U_PRG_HS_ZERO = "0b000000";
	parameter U_PRG_RXHS_SETTLE = "0b000000";
	parameter UC_PRG_HS_PREPARE = "1P0_TXCLKESC";
	parameter UC_PRG_HS_TRAIL = "0b00000";
	parameter UC_PRG_HS_ZERO = "0b0000000";
	parameter UC_PRG_RXHS_SETTLE = "0b000000";

endmodule

module DQSBUF_CORE (BTDETECT, BURSTDETECT, DATAVALID, DQSI, DQSW, DQSWRD, PAUSE, RDCLKSEL3, RDCLKSEL2, RDCLKSEL1, RDCLKSEL0, RDDIR, RDLOADN, RDPNTR2, RDPNTR1, RDPNTR0, READ3, READ2, READ1, READ0, READCOUT, READMOVE, RST, SCLK, SELCLK, DQSR90, DQSW270, WRCOUT, WRDIR, WRLOAD_N, WRLVCOUT, WRLVDIR, WRLVLOAD_N, WRLVMOVE, WRMOVE, WRPNTR2, WRPNTR1, WRPNTR0, ECLKIN, RSTSMCNT, DLLCODE8, DLLCODE7, DLLCODE6, DLLCODE5, DLLCODE4, DLLCODE3, DLLCODE2, DLLCODE1, DLLCODE0); //synthesis syn_black_box syn_lib_cell=1

	output BTDETECT;
	output BURSTDETECT;
	output DATAVALID;
	input DQSI;
	output DQSW;
	output DQSWRD;
	input PAUSE;
	input RDCLKSEL3;
	input RDCLKSEL2;
	input RDCLKSEL1;
	input RDCLKSEL0;
	input RDDIR;
	input RDLOADN;
	output RDPNTR2;
	output RDPNTR1;
	output RDPNTR0;
	input READ3;
	input READ2;
	input READ1;
	input READ0;
	output READCOUT;
	input READMOVE;
	input RST;
	input SCLK;
	input SELCLK;
	output DQSR90;
	output DQSW270;
	output WRCOUT;
	input WRDIR;
	input WRLOAD_N;
	output WRLVCOUT;
	input WRLVDIR;
	input WRLVLOAD_N;
	input WRLVMOVE;
	input WRMOVE;
	output WRPNTR2;
	output WRPNTR1;
	output WRPNTR0;
	input ECLKIN;
	input RSTSMCNT;
	input DLLCODE8;
	input DLLCODE7;
	input DLLCODE6;
	input DLLCODE5;
	input DLLCODE4;
	input DLLCODE3;
	input DLLCODE2;
	input DLLCODE1;
	input DLLCODE0;

	parameter GSR = "ENABLED";
	parameter ENABLE_FIFO = "DISABLED";
	parameter FORCE_READ = "DISABLED";
	parameter FREE_WHEEL = "DDR";
	parameter MODX = "NOT_USED";
	parameter MT_EN_READ = "DISABLED";
	parameter MT_EN_WRITE = "DISABLED";
	parameter MT_EN_WRITE_LEVELING = "DISABLED";
	parameter RD_PNTR = "0b000";
	parameter READ_ENABLE = "DISABLED";
	parameter RX_CENTERED = "ENABLED";
	parameter S_READ = "0";
	parameter S_WRITE = "0";
	parameter SIGN_READ = "POSITIVE";
	parameter SIGN_WRITE = "POSITIVE";
	parameter UPDATE_QU = "UP1_AND_UP0_SAME";
	parameter WRITE_ENABLE = "DISABLED";
	parameter SEL_READ_BIT_ENABLE_CYCLES = "NORMAL";
	parameter BYPASS_WR_LEVEL_SMTH_LATCH = "SMOOTHING_PATH";
	parameter BYPASS_WR_SMTH_LATCH = "SMOOTHING_PATH";
	parameter BYPASS_READ_SMTH_LATCH = "SMOOTHING_PATH";

endmodule

module ECLKDIV_CORE (DIVOUT, DIVRST, ECLKIN, SLIP, TESTINP3, TESTINP2, TESTINP1, TESTINP0); //synthesis syn_black_box syn_lib_cell=1

	output DIVOUT;
	input DIVRST;
	input ECLKIN;
	input SLIP;
	input TESTINP3;
	input TESTINP2;
	input TESTINP1;
	input TESTINP0;

	parameter ECLK_DIV = "DISABLE";
	parameter GSR = "ENABLED";

endmodule

module ECLKSYNC_CORE (ECLKIN, ECLKOUT, STOP); //synthesis syn_black_box syn_lib_cell=1

	input ECLKIN;
	output ECLKOUT;
	input STOP;

	parameter STOP_EN = "DISABLE";

endmodule

module FBMUX_CORE (ENEXT, FBKCK, LGYRDYN, INTLOCK, WKUPSYNC, FBKCLK15, FBKCLK14, FBKCLK13, FBKCLK12, FBKCLK11, FBKCLK10, FBKCLK9, FBKCLK8, FBKCLK7, FBKCLK6, FBKCLK5, FBKCLK4, FBKCLK3, FBKCLK2, FBKCLK1, FBKCLK0); //synthesis syn_black_box syn_lib_cell=1

	output ENEXT;
	output FBKCK;
	input LGYRDYN;
	input INTLOCK;
	input WKUPSYNC;
	input FBKCLK15;
	input FBKCLK14;
	input FBKCLK13;
	input FBKCLK12;
	input FBKCLK11;
	input FBKCLK10;
	input FBKCLK9;
	input FBKCLK8;
	input FBKCLK7;
	input FBKCLK6;
	input FBKCLK5;
	input FBKCLK4;
	input FBKCLK3;
	input FBKCLK2;
	input FBKCLK1;
	input FBKCLK0;

	parameter INTFB = "IGNORED";
	parameter SEL_FBK = "DIVA";
	parameter CLKMUX_FB = "CMUX_CLKOP";
	parameter INTFBKDEL_SEL = "DISABLED";

endmodule

module I2CFIFO_CORE (ALTSCLIN, ALTSCLOEN, ALTSCLOUT, ALTSDAIN, ALTSDAOEN, ALTSDAOUT, BUSBUSY, FIFORESET, I2CLSRRSTN, INSLEEP, IRQ, LMMICLK, LMMIOFFSET5, LMMIOFFSET4, LMMIOFFSET3, LMMIOFFSET2, LMMIOFFSET1, LMMIOFFSET0, LMMIRDATA7, LMMIRDATA6, LMMIRDATA5, LMMIRDATA4, LMMIRDATA3, LMMIRDATA2, LMMIRDATA1, LMMIRDATA0, LMMIRDATAVALID, LMMIREADY, LMMIREQUEST, LMMIRESETN, LMMIWDATA7, LMMIWDATA6, LMMIWDATA5, LMMIWDATA4, LMMIWDATA3, LMMIWDATA2, LMMIWDATA1, LMMIWDATA0, LMMIWRRDN, MRDCMPL, OPCGLOADCLK, RXFIFOAF, RXFIFOE, RXFIFOF, SCANCLK, SCANRST, SCLIN, SCLOE, SCLOEN, SCLOUT, SDAIN, SDAOE, SDAOEN, SDAOUT, SLEEPCLKSELN, SLVADDRMATCH, SLVADDRMATCHSCL, SRDWR, TXFIFOAE, TXFIFOE, TXFIFOF); //synthesis syn_black_box syn_lib_cell=1

	input ALTSCLIN;
	output ALTSCLOEN;
	output ALTSCLOUT;
	input ALTSDAIN;
	output ALTSDAOEN;
	output ALTSDAOUT;
	output BUSBUSY;
	input FIFORESET;
	input I2CLSRRSTN;
	output INSLEEP;
	output IRQ;
	input LMMICLK;
	input LMMIOFFSET5;
	input LMMIOFFSET4;
	input LMMIOFFSET3;
	input LMMIOFFSET2;
	input LMMIOFFSET1;
	input LMMIOFFSET0;
	output LMMIRDATA7;
	output LMMIRDATA6;
	output LMMIRDATA5;
	output LMMIRDATA4;
	output LMMIRDATA3;
	output LMMIRDATA2;
	output LMMIRDATA1;
	output LMMIRDATA0;
	output LMMIRDATAVALID;
	output LMMIREADY;
	input LMMIREQUEST;
	input LMMIRESETN;
	input LMMIWDATA7;
	input LMMIWDATA6;
	input LMMIWDATA5;
	input LMMIWDATA4;
	input LMMIWDATA3;
	input LMMIWDATA2;
	input LMMIWDATA1;
	input LMMIWDATA0;
	input LMMIWRRDN;
	output MRDCMPL;
	input OPCGLOADCLK;
	output RXFIFOAF;
	output RXFIFOE;
	output RXFIFOF;
	input SCANCLK;
	input SCANRST;
	input SCLIN;
	output SCLOE;
	output SCLOEN;
	output SCLOUT;
	input SDAIN;
	output SDAOE;
	output SDAOEN;
	output SDAOUT;
	input SLEEPCLKSELN;
	output SLVADDRMATCH;
	output SLVADDRMATCHSCL;
	output SRDWR;
	output TXFIFOAE;
	output TXFIFOE;
	output TXFIFOF;

	parameter BRNBASEDELAY = "0b0000";
	parameter CR1CKDIS = "EN";
	parameter CR1FIFOMODE = "REG";
	parameter CR1GCEN = "DIS";
	parameter CR1I2CEN = "DIS";
	parameter CR1SDADELSEL = "NDLY0";
	parameter CR1SLPCLKEN = "DIS";
	parameter CR2CORERSTN = "DIS";
	parameter CR2HARDTIE = "TIE";
	parameter CR2INTCLREN = "DIS";
	parameter CR2MRDCMPLWKUP = "DIS";
	parameter CR2RXFIFOAFWKUP = "DIS";
	parameter CR2SLVADDRWKUP = "DIS";
	parameter GSR = "ENABLED";
    parameter I2CADDRSEL = "7BIT";
	parameter I2CRXFIFOAFVAL = "0b00000";
	parameter I2CSLVADDRA = "0b0000000000";
	parameter I2CTXFIFOAEVAL = "0b0000";
	parameter INTARBLIE = "DIS";
	parameter INTBUSFREEIE = "DIS";
	parameter INTHGCIE = "DIS";
	parameter INTMRDCMPLIE = "DIS";
	parameter INTRNACKIEORRSVD = "DIS";
	parameter INTRSVDORTROEIE = "DIS";
	parameter INTRSVDORTRRDYIE = "DIS";
	parameter INTRXOVERFIEORRSVD = "DIS";
	parameter INTRXUNDERFIE = "DIS";
	parameter INTTXOVERFIE = "DIS";
	parameter INTTXSERRIEORRSVD = "DIS";
	parameter LMMI_EXTRA_ONE = "DIS";
	parameter LMMI_EXTRA_TWO = "DIS";
	parameter NCRALTIOEN = "FABRIC";
	parameter NCRFILTERDIS = "EN";
	parameter NCRSDAINDLYEN = "DIS";
	parameter NCRSDAOUTDLYEN = "DIS";
	parameter NONUSRTESTSOFTTRIMEN = "DIS";
	parameter NONUSRTSTSOFTTRIMVALUE = "0b000";
	parameter REGI2CBR = "0b0000000000";
	parameter TSPTIMERVALUE = "0b10010010111";

endmodule

module LRAM_CORE (ADA13, ADA12, ADA11, ADA10, ADA9, ADA8, ADA7, ADA6, ADA5, ADA4, ADA3, ADA2, ADA1, ADA0, ADB13, ADB12, ADB11, ADB10, ADB9, ADB8, ADB7, ADB6, ADB5, ADB4, ADB3, ADB2, ADB1, ADB0, BENA_N3, BENA_N2, BENA_N1, BENA_N0, BENB_N3, BENB_N2, BENB_N1, BENB_N0, CEA, CEB, CLK, CSA, CSB, DIA31, DIA30, DIA29, DIA28, DIA27, DIA26, DIA25, DIA24, DIA23, DIA22, DIA21, DIA20, DIA19, DIA18, DIA17, DIA16, DIA15, DIA14, DIA13, DIA12, DIA11, DIA10, DIA9, DIA8, DIA7, DIA6, DIA5, DIA4, DIA3, DIA2, DIA1, DIA0, DIB31, DIB30, DIB29, DIB28, DIB27, DIB26, DIB25, DIB24, DIB23, DIB22, DIB21, DIB20, DIB19, DIB18, DIB17, DIB16, DIB15, DIB14, DIB13, DIB12, DIB11, DIB10, DIB9, DIB8, DIB7, DIB6, DIB5, DIB4, DIB3, DIB2, DIB1, DIB0, DOA31, DOA30, DOA29, DOA28, DOA27, DOA26, DOA25, DOA24, DOA23, DOA22, DOA21, DOA20, DOA19, DOA18, DOA17, DOA16, DOA15, DOA14, DOA13, DOA12, DOA11, DOA10, DOA9, DOA8, DOA7, DOA6, DOA5, DOA4, DOA3, DOA2, DOA1, DOA0, DOB31, DOB30, DOB29, DOB28, DOB27, DOB26, DOB25, DOB24, DOB23, DOB22, DOB21, DOB20, DOB19, DOB18, DOB17, DOB16, DOB15, DOB14, DOB13, DOB12, DOB11, DOB10, DOB9, DOB8, DOB7, DOB6, DOB5, DOB4, DOB3, DOB2, DOB1, DOB0, DPS, ERRDECA1, ERRDECA0, ERRDECB1, ERRDECB0, IGN, INITN, OCEA, OCEB, OEA, OEB, RSTA, RSTB, STDBYN, TBISTN, WEA, WEB, ERRDET, LRAMREADY, OPCGLOADCLK, SCANCLK, SCANRST); //synthesis syn_black_box syn_lib_cell=1

	input ADA13;
	input ADA12;
	input ADA11;
	input ADA10;
	input ADA9;
	input ADA8;
	input ADA7;
	input ADA6;
	input ADA5;
	input ADA4;
	input ADA3;
	input ADA2;
	input ADA1;
	input ADA0;
	input ADB13;
	input ADB12;
	input ADB11;
	input ADB10;
	input ADB9;
	input ADB8;
	input ADB7;
	input ADB6;
	input ADB5;
	input ADB4;
	input ADB3;
	input ADB2;
	input ADB1;
	input ADB0;
	input BENA_N3;
	input BENA_N2;
	input BENA_N1;
	input BENA_N0;
	input BENB_N3;
	input BENB_N2;
	input BENB_N1;
	input BENB_N0;
	input CEA;
	input CEB;
	input CLK;
	input CSA;
	input CSB;
	input DIA31;
	input DIA30;
	input DIA29;
	input DIA28;
	input DIA27;
	input DIA26;
	input DIA25;
	input DIA24;
	input DIA23;
	input DIA22;
	input DIA21;
	input DIA20;
	input DIA19;
	input DIA18;
	input DIA17;
	input DIA16;
	input DIA15;
	input DIA14;
	input DIA13;
	input DIA12;
	input DIA11;
	input DIA10;
	input DIA9;
	input DIA8;
	input DIA7;
	input DIA6;
	input DIA5;
	input DIA4;
	input DIA3;
	input DIA2;
	input DIA1;
	input DIA0;
	input DIB31;
	input DIB30;
	input DIB29;
	input DIB28;
	input DIB27;
	input DIB26;
	input DIB25;
	input DIB24;
	input DIB23;
	input DIB22;
	input DIB21;
	input DIB20;
	input DIB19;
	input DIB18;
	input DIB17;
	input DIB16;
	input DIB15;
	input DIB14;
	input DIB13;
	input DIB12;
	input DIB11;
	input DIB10;
	input DIB9;
	input DIB8;
	input DIB7;
	input DIB6;
	input DIB5;
	input DIB4;
	input DIB3;
	input DIB2;
	input DIB1;
	input DIB0;
	output DOA31;
	output DOA30;
	output DOA29;
	output DOA28;
	output DOA27;
	output DOA26;
	output DOA25;
	output DOA24;
	output DOA23;
	output DOA22;
	output DOA21;
	output DOA20;
	output DOA19;
	output DOA18;
	output DOA17;
	output DOA16;
	output DOA15;
	output DOA14;
	output DOA13;
	output DOA12;
	output DOA11;
	output DOA10;
	output DOA9;
	output DOA8;
	output DOA7;
	output DOA6;
	output DOA5;
	output DOA4;
	output DOA3;
	output DOA2;
	output DOA1;
	output DOA0;
	output DOB31;
	output DOB30;
	output DOB29;
	output DOB28;
	output DOB27;
	output DOB26;
	output DOB25;
	output DOB24;
	output DOB23;
	output DOB22;
	output DOB21;
	output DOB20;
	output DOB19;
	output DOB18;
	output DOB17;
	output DOB16;
	output DOB15;
	output DOB14;
	output DOB13;
	output DOB12;
	output DOB11;
	output DOB10;
	output DOB9;
	output DOB8;
	output DOB7;
	output DOB6;
	output DOB5;
	output DOB4;
	output DOB3;
	output DOB2;
	output DOB1;
	output DOB0;
	input DPS;
	output ERRDECA1;
	output ERRDECA0;
	output ERRDECB1;
	output ERRDECB0;
	input IGN;
	input INITN;
	input OCEA;
	input OCEB;
	output OEA;
	output OEB;
	input RSTA;
	input RSTB;
	input STDBYN;
	input TBISTN;
	input WEA;
	input WEB;
	output ERRDET;
	output LRAMREADY;
	input OPCGLOADCLK;
	input SCANCLK;
	input SCANRST;

	parameter INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_40 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_41 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_42 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_43 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_44 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_45 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_46 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_47 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_48 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_49 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_4A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_4B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_4C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_4D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_4E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_4F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_50 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_51 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_52 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_53 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_54 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_55 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_56 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_57 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_58 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_59 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_5A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_5B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_5C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_5D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_5E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_5F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_60 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_61 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_62 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_63 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_64 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_65 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_66 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_67 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_68 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_69 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_6A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_6B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_6C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_6D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_6E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_6F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_70 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_71 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_72 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_73 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_74 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_75 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_76 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_77 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_78 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_79 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_7A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_7B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_7C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_7D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_7E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_7F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter ASYNC_RST_RELEASE = "SYNC";
	parameter CFG_INIT_ID = "0b00000000000";
	parameter DATA_PRESERVE = "DISABLE";
	parameter EBR_SP_EN = "DISABLE";
	parameter ECC_BYTE_SEL = "ECC_EN";
	parameter GSR = "ENABLED";
	parameter OUT_REGMODE_A = "NO_REG";
	parameter OUT_REGMODE_B = "NO_REG";
	parameter RESETMODE = "SYNC";
	parameter RST_AB_EN = "RESET_AB_DISABLE";
	parameter SP_EN = "DISABLE";
	parameter UNALIGNED_READ = "DISABLE";

endmodule

module MULT18_CORE (SFTCTRL3, SFTCTRL2, SFTCTRL1, SFTCTRL0, ARHSIGN, BRHSIGN, ARH8, ARH7, ARH6, ARH5, ARH4, ARH3, ARH2, ARH1, ARH0, BRH8, BRH7, BRH6, BRH5, BRH4, BRH3, BRH2, BRH1, BRH0, ARL8, ARL7, ARL6, ARL5, ARL4, ARL3, ARL2, ARL1, ARL0, BRL8, BRL7, BRL6, BRL5, BRL4, BRL3, BRL2, BRL1, BRL0, PL1819, PL1818, PL1817, PL1816, PL1815, PL1814, PL1813, PL1812, PL1811, PL1810, PL189, PL188, PL187, PL186, PL185, PL184, PL183, PL182, PL181, PL180, PH1819, PH1818, PH1817, PH1816, PH1815, PH1814, PH1813, PH1812, PH1811, PH1810, PH189, PH188, PH187, PH186, PH185, PH184, PH183, PH182, PH181, PH180, SIGNED18, P3637, P3636, P3635, P3634, P3633, P3632, P3631, P3630, P3629, P3628, P3627, P3626, P3625, P3624, P3623, P3622, P3621, P3620, P3619, P3618, P3617, P3616, P3615, P3614, P3613, P3612, P3611, P3610, P369, P368, P367, P366, P365, P364, P363, P362, P361, P360, ROUNDEN); //synthesis syn_black_box syn_lib_cell=1

	input SFTCTRL3;
	input SFTCTRL2;
	input SFTCTRL1;
	input SFTCTRL0;
	input ARHSIGN;
	input BRHSIGN;
	input ARH8;
	input ARH7;
	input ARH6;
	input ARH5;
	input ARH4;
	input ARH3;
	input ARH2;
	input ARH1;
	input ARH0;
	input BRH8;
	input BRH7;
	input BRH6;
	input BRH5;
	input BRH4;
	input BRH3;
	input BRH2;
	input BRH1;
	input BRH0;
	input ARL8;
	input ARL7;
	input ARL6;
	input ARL5;
	input ARL4;
	input ARL3;
	input ARL2;
	input ARL1;
	input ARL0;
	input BRL8;
	input BRL7;
	input BRL6;
	input BRL5;
	input BRL4;
	input BRL3;
	input BRL2;
	input BRL1;
	input BRL0;
	input PL1819;
	input PL1818;
	input PL1817;
	input PL1816;
	input PL1815;
	input PL1814;
	input PL1813;
	input PL1812;
	input PL1811;
	input PL1810;
	input PL189;
	input PL188;
	input PL187;
	input PL186;
	input PL185;
	input PL184;
	input PL183;
	input PL182;
	input PL181;
	input PL180;
	input PH1819;
	input PH1818;
	input PH1817;
	input PH1816;
	input PH1815;
	input PH1814;
	input PH1813;
	input PH1812;
	input PH1811;
	input PH1810;
	input PH189;
	input PH188;
	input PH187;
	input PH186;
	input PH185;
	input PH184;
	input PH183;
	input PH182;
	input PH181;
	input PH180;
	output SIGNED18;
	output P3637;
	output P3636;
	output P3635;
	output P3634;
	output P3633;
	output P3632;
	output P3631;
	output P3630;
	output P3629;
	output P3628;
	output P3627;
	output P3626;
	output P3625;
	output P3624;
	output P3623;
	output P3622;
	output P3621;
	output P3620;
	output P3619;
	output P3618;
	output P3617;
	output P3616;
	output P3615;
	output P3614;
	output P3613;
	output P3612;
	output P3611;
	output P3610;
	output P369;
	output P368;
	output P367;
	output P366;
	output P365;
	output P364;
	output P363;
	output P362;
	output P361;
	output P360;
	input ROUNDEN;

	parameter SFTEN = "DISABLED";
	parameter MULT18X18 = "ENABLED";
	parameter ROUNDHALFUP = "DISABLED";
	parameter ROUNDRTZI = "ROUND_TO_ZERO";
	parameter ROUNDBIT = "ROUND_TO_BIT0";

endmodule

module MULT18X36_CORE (SFTCTRL3, SFTCTRL2, SFTCTRL1, SFTCTRL0, PH3637, PH3636, PH3635, PH3634, PH3633, PH3632, PH3631, PH3630, PH3629, PH3628, PH3627, PH3626, PH3625, PH3624, PH3623, PH3622, PH3621, PH3620, PH3619, PH3618, PH3617, PH3616, PH3615, PH3614, PH3613, PH3612, PH3611, PH3610, PH369, PH368, PH367, PH366, PH365, PH364, PH363, PH362, PH361, PH360, PL3637, PL3636, PL3635, PL3634, PL3633, PL3632, PL3631, PL3630, PL3629, PL3628, PL3627, PL3626, PL3625, PL3624, PL3623, PL3622, PL3621, PL3620, PL3619, PL3618, PL3617, PL3616, PL3615, PL3614, PL3613, PL3612, PL3611, PL3610, PL369, PL368, PL367, PL366, PL365, PL364, PL363, PL362, PL361, PL360, SGNED18H, SGNED18L, P7272, P7271, P7270, P7269, P7268, P7267, P7266, P7265, P7264, P7263, P7262, P7261, P7260, P7259, P7258, P7257, P7256, P7255, P7254, P7253, P7252, P7251, P7250, P7249, P7248, P7247, P7246, P7245, P7244, P7243, P7242, P7241, P7240, P7239, P7238, P7237, P7236, P7235, P7234, P7233, P7232, P7231, P7230, P7229, P7228, P7227, P7226, P7225, P7224, P7223, P7222, P7221, P7220, P7219, P7218, P7217, P7216, P7215, P7214, P7213, P7212, P7211, P7210, P729, P728, P727, P726, P725, P724, P723, P722, P721, P720, ROUNDEN); //synthesis syn_black_box syn_lib_cell=1

	input SFTCTRL3;
	input SFTCTRL2;
	input SFTCTRL1;
	input SFTCTRL0;
	input PH3637;
	input PH3636;
	input PH3635;
	input PH3634;
	input PH3633;
	input PH3632;
	input PH3631;
	input PH3630;
	input PH3629;
	input PH3628;
	input PH3627;
	input PH3626;
	input PH3625;
	input PH3624;
	input PH3623;
	input PH3622;
	input PH3621;
	input PH3620;
	input PH3619;
	input PH3618;
	input PH3617;
	input PH3616;
	input PH3615;
	input PH3614;
	input PH3613;
	input PH3612;
	input PH3611;
	input PH3610;
	input PH369;
	input PH368;
	input PH367;
	input PH366;
	input PH365;
	input PH364;
	input PH363;
	input PH362;
	input PH361;
	input PH360;
	input PL3637;
	input PL3636;
	input PL3635;
	input PL3634;
	input PL3633;
	input PL3632;
	input PL3631;
	input PL3630;
	input PL3629;
	input PL3628;
	input PL3627;
	input PL3626;
	input PL3625;
	input PL3624;
	input PL3623;
	input PL3622;
	input PL3621;
	input PL3620;
	input PL3619;
	input PL3618;
	input PL3617;
	input PL3616;
	input PL3615;
	input PL3614;
	input PL3613;
	input PL3612;
	input PL3611;
	input PL3610;
	input PL369;
	input PL368;
	input PL367;
	input PL366;
	input PL365;
	input PL364;
	input PL363;
	input PL362;
	input PL361;
	input PL360;
	input SGNED18H;
	input SGNED18L;
	output P7272;
	output P7271;
	output P7270;
	output P7269;
	output P7268;
	output P7267;
	output P7266;
	output P7265;
	output P7264;
	output P7263;
	output P7262;
	output P7261;
	output P7260;
	output P7259;
	output P7258;
	output P7257;
	output P7256;
	output P7255;
	output P7254;
	output P7253;
	output P7252;
	output P7251;
	output P7250;
	output P7249;
	output P7248;
	output P7247;
	output P7246;
	output P7245;
	output P7244;
	output P7243;
	output P7242;
	output P7241;
	output P7240;
	output P7239;
	output P7238;
	output P7237;
	output P7236;
	output P7235;
	output P7234;
	output P7233;
	output P7232;
	output P7231;
	output P7230;
	output P7229;
	output P7228;
	output P7227;
	output P7226;
	output P7225;
	output P7224;
	output P7223;
	output P7222;
	output P7221;
	output P7220;
	output P7219;
	output P7218;
	output P7217;
	output P7216;
	output P7215;
	output P7214;
	output P7213;
	output P7212;
	output P7211;
	output P7210;
	output P729;
	output P728;
	output P727;
	output P726;
	output P725;
	output P724;
	output P723;
	output P722;
	output P721;
	output P720;
	input ROUNDEN;

	parameter SFTEN = "DISABLED";
	parameter MULT18X36 = "ENABLED";
	parameter MULT36 = "DISABLED";
	parameter MULT36X36H = "USED_AS_LOWER_BIT_GENERATION";
	parameter ROUNDHALFUP = "DISABLED";
	parameter ROUNDRTZI = "ROUND_TO_ZERO";
	parameter ROUNDBIT = "ROUND_TO_BIT0";

endmodule

module MULT36_CORE (PH7272, PH7271, PH7270, PH7269, PH7268, PH7267, PH7266, PH7265, PH7264, PH7263, PH7262, PH7261, PH7260, PH7259, PH7258, PH7257, PH7256, PH7255, PH7254, PH7253, PH7252, PH7251, PH7250, PH7249, PH7248, PH7247, PH7246, PH7245, PH7244, PH7243, PH7242, PH7241, PH7240, PH7239, PH7238, PH7237, PH7236, PH7235, PH7234, PH7233, PH7232, PH7231, PH7230, PH7229, PH7228, PH7227, PH7226, PH7225, PH7224, PH7223, PH7222, PH7221, PH7220, PH7219, PH7218, PH7217, PH7216, PH7215, PH7214, PH7213, PH7212, PH7211, PH7210, PH729, PH728, PH727, PH726, PH725, PH724, PH723, PH722, PH721, PH720, PL7272, PL7271, PL7270, PL7269, PL7268, PL7267, PL7266, PL7265, PL7264, PL7263, PL7262, PL7261, PL7260, PL7259, PL7258, PL7257, PL7256, PL7255, PL7254, PL7253, PL7252, PL7251, PL7250, PL7249, PL7248, PL7247, PL7246, PL7245, PL7244, PL7243, PL7242, PL7241, PL7240, PL7239, PL7238, PL7237, PL7236, PL7235, PL7234, PL7233, PL7232, PL7231, PL7230, PL7229, PL7228, PL7227, PL7226, PL7225, PL7224, PL7223, PL7222, PL7221, PL7220, PL7219, PL7218, PL7217, PL7216, PL7215, PL7214, PL7213, PL7212, PL7211, PL7210, PL729, PL728, PL727, PL726, PL725, PL724, PL723, PL722, PL721, PL720, PML7271, PML7270, PML7269, PML7268, PML7267, PML7266, PML7265, PML7264, PML7263, PML7262, PML7261, PML7260, PML7259, PML7258, PML7257, PML7256, PML7255, PML7254, PML7253, PML7252, PML7251, PML7250, PML7249, PML7248, PML7247, PML7246, PML7245, PML7244, PML7243, PML7242, PML7241, PML7240, PML7239, PML7238, PML7237, PML7236, PML7235, PML7234, PML7233, PML7232, PML7231, PML7230, PML7229, PML7228, PML7227, PML7226, PML7225, PML7224, PML7223, PML7222, PML7221, PML7220, PML7219, PML7218, PML7217, PML7216, PML7215, PML7214, PML7213, PML7212, PML7211, PML7210, PML729, PML728, PML727, PML726, PML725, PML724, PML723, PML722, PML721, PML720, PMH7271, PMH7270, PMH7269, PMH7268, PMH7267, PMH7266, PMH7265, PMH7264, PMH7263, PMH7262, PMH7261, PMH7260, PMH7259, PMH7258, PMH7257, PMH7256, PMH7255, PMH7254, PMH7253, PMH7252, PMH7251, PMH7250, PMH7249, PMH7248, PMH7247, PMH7246, PMH7245, PMH7244, PMH7243, PMH7242, PMH7241, PMH7240, PMH7239, PMH7238, PMH7237, PMH7236, PMH7235, PMH7234, PMH7233, PMH7232, PMH7231, PMH7230, PMH7229, PMH7228, PMH7227, PMH7226, PMH7225, PMH7224, PMH7223, PMH7222, PMH7221, PMH7220, PMH7219, PMH7218, PMH7217, PMH7216, PMH7215, PMH7214, PMH7213, PMH7212, PMH7211, PMH7210, PMH729, PMH728, PMH727, PMH726, PMH725, PMH724, PMH723, PMH722, PMH721, PMH720); //synthesis syn_black_box syn_lib_cell=1

	input PH7272;
	input PH7271;
	input PH7270;
	input PH7269;
	input PH7268;
	input PH7267;
	input PH7266;
	input PH7265;
	input PH7264;
	input PH7263;
	input PH7262;
	input PH7261;
	input PH7260;
	input PH7259;
	input PH7258;
	input PH7257;
	input PH7256;
	input PH7255;
	input PH7254;
	input PH7253;
	input PH7252;
	input PH7251;
	input PH7250;
	input PH7249;
	input PH7248;
	input PH7247;
	input PH7246;
	input PH7245;
	input PH7244;
	input PH7243;
	input PH7242;
	input PH7241;
	input PH7240;
	input PH7239;
	input PH7238;
	input PH7237;
	input PH7236;
	input PH7235;
	input PH7234;
	input PH7233;
	input PH7232;
	input PH7231;
	input PH7230;
	input PH7229;
	input PH7228;
	input PH7227;
	input PH7226;
	input PH7225;
	input PH7224;
	input PH7223;
	input PH7222;
	input PH7221;
	input PH7220;
	input PH7219;
	input PH7218;
	input PH7217;
	input PH7216;
	input PH7215;
	input PH7214;
	input PH7213;
	input PH7212;
	input PH7211;
	input PH7210;
	input PH729;
	input PH728;
	input PH727;
	input PH726;
	input PH725;
	input PH724;
	input PH723;
	input PH722;
	input PH721;
	input PH720;
	input PL7272;
	input PL7271;
	input PL7270;
	input PL7269;
	input PL7268;
	input PL7267;
	input PL7266;
	input PL7265;
	input PL7264;
	input PL7263;
	input PL7262;
	input PL7261;
	input PL7260;
	input PL7259;
	input PL7258;
	input PL7257;
	input PL7256;
	input PL7255;
	input PL7254;
	input PL7253;
	input PL7252;
	input PL7251;
	input PL7250;
	input PL7249;
	input PL7248;
	input PL7247;
	input PL7246;
	input PL7245;
	input PL7244;
	input PL7243;
	input PL7242;
	input PL7241;
	input PL7240;
	input PL7239;
	input PL7238;
	input PL7237;
	input PL7236;
	input PL7235;
	input PL7234;
	input PL7233;
	input PL7232;
	input PL7231;
	input PL7230;
	input PL7229;
	input PL7228;
	input PL7227;
	input PL7226;
	input PL7225;
	input PL7224;
	input PL7223;
	input PL7222;
	input PL7221;
	input PL7220;
	input PL7219;
	input PL7218;
	input PL7217;
	input PL7216;
	input PL7215;
	input PL7214;
	input PL7213;
	input PL7212;
	input PL7211;
	input PL7210;
	input PL729;
	input PL728;
	input PL727;
	input PL726;
	input PL725;
	input PL724;
	input PL723;
	input PL722;
	input PL721;
	input PL720;
	output PML7271;
	output PML7270;
	output PML7269;
	output PML7268;
	output PML7267;
	output PML7266;
	output PML7265;
	output PML7264;
	output PML7263;
	output PML7262;
	output PML7261;
	output PML7260;
	output PML7259;
	output PML7258;
	output PML7257;
	output PML7256;
	output PML7255;
	output PML7254;
	output PML7253;
	output PML7252;
	output PML7251;
	output PML7250;
	output PML7249;
	output PML7248;
	output PML7247;
	output PML7246;
	output PML7245;
	output PML7244;
	output PML7243;
	output PML7242;
	output PML7241;
	output PML7240;
	output PML7239;
	output PML7238;
	output PML7237;
	output PML7236;
	output PML7235;
	output PML7234;
	output PML7233;
	output PML7232;
	output PML7231;
	output PML7230;
	output PML7229;
	output PML7228;
	output PML7227;
	output PML7226;
	output PML7225;
	output PML7224;
	output PML7223;
	output PML7222;
	output PML7221;
	output PML7220;
	output PML7219;
	output PML7218;
	output PML7217;
	output PML7216;
	output PML7215;
	output PML7214;
	output PML7213;
	output PML7212;
	output PML7211;
	output PML7210;
	output PML729;
	output PML728;
	output PML727;
	output PML726;
	output PML725;
	output PML724;
	output PML723;
	output PML722;
	output PML721;
	output PML720;
	output PMH7271;
	output PMH7270;
	output PMH7269;
	output PMH7268;
	output PMH7267;
	output PMH7266;
	output PMH7265;
	output PMH7264;
	output PMH7263;
	output PMH7262;
	output PMH7261;
	output PMH7260;
	output PMH7259;
	output PMH7258;
	output PMH7257;
	output PMH7256;
	output PMH7255;
	output PMH7254;
	output PMH7253;
	output PMH7252;
	output PMH7251;
	output PMH7250;
	output PMH7249;
	output PMH7248;
	output PMH7247;
	output PMH7246;
	output PMH7245;
	output PMH7244;
	output PMH7243;
	output PMH7242;
	output PMH7241;
	output PMH7240;
	output PMH7239;
	output PMH7238;
	output PMH7237;
	output PMH7236;
	output PMH7235;
	output PMH7234;
	output PMH7233;
	output PMH7232;
	output PMH7231;
	output PMH7230;
	output PMH7229;
	output PMH7228;
	output PMH7227;
	output PMH7226;
	output PMH7225;
	output PMH7224;
	output PMH7223;
	output PMH7222;
	output PMH7221;
	output PMH7220;
	output PMH7219;
	output PMH7218;
	output PMH7217;
	output PMH7216;
	output PMH7215;
	output PMH7214;
	output PMH7213;
	output PMH7212;
	output PMH7211;
	output PMH7210;
	output PMH729;
	output PMH728;
	output PMH727;
	output PMH726;
	output PMH725;
	output PMH724;
	output PMH723;
	output PMH722;
	output PMH721;
	output PMH720;

	parameter MULT36X36 = "ENABLED";

endmodule

module MULT9_CORE (A8, A7, A6, A5, A4, A3, A2, A1, A0, ASIGNED, BR8, BR7, BR6, BR5, BR4, BR3, BR2, BR1, BR0, AS18, AS17, AS16, AS15, AS14, AS13, AS12, AS11, AS10, AS28, AS27, AS26, AS25, AS24, AS23, AS22, AS21, AS20, ASSIGNED1, ASSIGNED2, BRSIGNED, CLK, CEA, RSTA, AO8, AO7, AO6, AO5, AO4, AO3, AO2, AO1, AO0, BO8, BO7, BO6, BO5, BO4, BO3, BO2, BO1, BO0, AOSIGNED, BOSIGNED, AR8, AR7, AR6, AR5, AR4, AR3, AR2, AR1, AR0, ARSIGNED, P1819, P1818, P1817, P1816, P1815, P1814, P1813, P1812, P1811, P1810, P189, P188, P187, P186, P185, P184, P183, P182, P181, P180, CEP, RSTP); //synthesis syn_black_box syn_lib_cell=1

	input A8;
	input A7;
	input A6;
	input A5;
	input A4;
	input A3;
	input A2;
	input A1;
	input A0;
	input ASIGNED;
	input BR8;
	input BR7;
	input BR6;
	input BR5;
	input BR4;
	input BR3;
	input BR2;
	input BR1;
	input BR0;
	input AS18;
	input AS17;
	input AS16;
	input AS15;
	input AS14;
	input AS13;
	input AS12;
	input AS11;
	input AS10;
	input AS28;
	input AS27;
	input AS26;
	input AS25;
	input AS24;
	input AS23;
	input AS22;
	input AS21;
	input AS20;
	input ASSIGNED1;
	input ASSIGNED2;
	input BRSIGNED;
	input CLK;
	input CEA;
	input RSTA;
	output AO8;
	output AO7;
	output AO6;
	output AO5;
	output AO4;
	output AO3;
	output AO2;
	output AO1;
	output AO0;
	output BO8;
	output BO7;
	output BO6;
	output BO5;
	output BO4;
	output BO3;
	output BO2;
	output BO1;
	output BO0;
	output AOSIGNED;
	output BOSIGNED;
	output AR8;
	output AR7;
	output AR6;
	output AR5;
	output AR4;
	output AR3;
	output AR2;
	output AR1;
	output AR0;
	output ARSIGNED;
	output P1819;
	output P1818;
	output P1817;
	output P1816;
	output P1815;
	output P1814;
	output P1813;
	output P1812;
	output P1811;
	output P1810;
	output P189;
	output P188;
	output P187;
	output P186;
	output P185;
	output P184;
	output P183;
	output P182;
	output P181;
	output P180;
	input CEP;
	input RSTP;

	parameter SIGNEDSTATIC_EN = "DISABLED";
	parameter ASIGNED_OPERAND_EN = "DISABLED";
	parameter BYPASS_MULT9 = "USED";
	parameter REGBYPSB = "REGISTER";
	parameter REGBYPSA1 = "REGISTER";
	parameter REGBYPSA2 = "REGISTER";
	parameter SHIFTA = "DISABLED";
	parameter SR_18BITSHIFT_EN = "DISABLED";
	parameter GSR = "ENABLED";
	parameter RESET = "SYNC";

endmodule

module OSC_CORE (HFCLKOUT, HFOUTEN, HFSDSCEN, HFTRMFAB8, HFTRMFAB7, HFTRMFAB6, HFTRMFAB5, HFTRMFAB4, HFTRMFAB3, HFTRMFAB2, HFTRMFAB1, HFTRMFAB0, LFCLKOUT, LFTRMFAB8, LFTRMFAB7, LFTRMFAB6, LFTRMFAB5, LFTRMFAB4, LFTRMFAB3, LFTRMFAB2, LFTRMFAB1, LFTRMFAB0, HFCLKCFG, HFSDCOUT); //synthesis syn_black_box syn_lib_cell=1

	output HFCLKOUT;
	input HFOUTEN;
	input HFSDSCEN;
	input HFTRMFAB8;
	input HFTRMFAB7;
	input HFTRMFAB6;
	input HFTRMFAB5;
	input HFTRMFAB4;
	input HFTRMFAB3;
	input HFTRMFAB2;
	input HFTRMFAB1;
	input HFTRMFAB0;
	output LFCLKOUT;
	input LFTRMFAB8;
	input LFTRMFAB7;
	input LFTRMFAB6;
	input LFTRMFAB5;
	input LFTRMFAB4;
	input LFTRMFAB3;
	input LFTRMFAB2;
	input LFTRMFAB1;
	input LFTRMFAB0;
	output HFCLKCFG;
	output HFSDCOUT;

	parameter DTR_EN = "ENABLED";
	parameter HF_CLK_DIV = "1";
	parameter HF_SED_SEC_DIV = "1";
	parameter HF_FABRIC_EN = "DISABLED";
	parameter HF_OSC_EN = "ENABLED";
	parameter HFDIV_FABRIC_EN = "ENABLED";
	parameter LF_FABRIC_EN = "DISABLED";
	parameter LF_OUTPUT_EN = "DISABLED";
	parameter DEBUG_N = "DISABLED";

endmodule

module PCIE_CORE (ACTACMD, ACTDR11, ACTEN, ACTHIGHZ, ACTMD, ACJNOUT, ACJPOUT, AUXCK, CKUSRI, CKUSRO, ECKIN, ECKIND2, ECKINDO, ERSTN, ERSTND2, ERXCKD2, ERXCKDO, ERXRSND2, ETXCKD2, ETXCKDO, ETXRSND2, FLR3, FLR2, FLR1, FLR0, FLRACK3, FLRACK2, FLRACK1, FLRACK0, MINTLEG3, MINTLEG2, MINTLEG1, MINTLEG0, MINTO, PERSTN, PMCTRL4, PMCTRL3, PMCTRL2, PMCTRL1, PMCTRL0, PMCTRLEN, PMDPAST4, PMDPAST3, PMDPAST2, PMDPAST1, PMDPAST0, PRMSGSD, PRNOSNP12, PRNOSNP11, PRNOSNP10, PRNOSNP9, PRNOSNP8, PRNOSNP7, PRNOSNP6, PRNOSNP5, PRNOSNP4, PRNOSNP3, PRNOSNP2, PRNOSNP1, PRNOSNP0, PRNSNPRE, PRSNOOP12, PRSNOOP11, PRSNOOP10, PRSNOOP9, PRSNOOP8, PRSNOOP7, PRSNOOP6, PRSNOOP5, PRSNOOP4, PRSNOOP3, PRSNOOP2, PRSNOOP1, PRSNOOP0, PRSNPRE, PPBDREG31, PPBDREG30, PPBDREG29, PPBDREG28, PPBDREG27, PPBDREG26, PPBDREG25, PPBDREG24, PPBDREG23, PPBDREG22, PPBDREG21, PPBDREG20, PPBDREG19, PPBDREG18, PPBDREG17, PPBDREG16, PPBDREG15, PPBDREG14, PPBDREG13, PPBDREG12, PPBDREG11, PPBDREG10, PPBDREG9, PPBDREG8, PPBDREG7, PPBDREG6, PPBDREG5, PPBDREG4, PPBDREG3, PPBDREG2, PPBDREG1, PPBDREG0, PPBDSEL7, PPBDSEL6, PPBDSEL5, PPBDSEL4, PPBDSEL3, PPBDSEL2, PPBDSEL1, PPBDSEL0, REXTCK, REXTRST, RSTUSRN, UDLLKUP, ULTSDIS, UPLLKUP, UTLLKUP, UCFGADDR11, UCFGADDR10, UCFGADDR9, UCFGADDR8, UCFGADDR7, UCFGADDR6, UCFGADDR5, UCFGADDR4, UCFGADDR3, UCFGADDR2, UCFGF2, UCFGF1, UCFGF0, UCFGRDD31, UCFGRDD30, UCFGRDD29, UCFGRDD28, UCFGRDD27, UCFGRDD26, UCFGRDD25, UCFGRDD24, UCFGRDD23, UCFGRDD22, UCFGRDD21, UCFGRDD20, UCFGRDD19, UCFGRDD18, UCFGRDD17, UCFGRDD16, UCFGRDD15, UCFGRDD14, UCFGRDD13, UCFGRDD12, UCFGRDD11, UCFGRDD10, UCFGRDD9, UCFGRDD8, UCFGRDD7, UCFGRDD6, UCFGRDD5, UCFGRDD4, UCFGRDD3, UCFGRDD2, UCFGRDD1, UCFGRDD0, UCFGRDE, UCFGRDY, UCFGSERD, UCFGVD, UCFGWRBE3, UCFGWRBE2, UCFGWRBE1, UCFGWRBE0, UCFGWRD31, UCFGWRD30, UCFGWRD29, UCFGWRD28, UCFGWRD27, UCFGWRD26, UCFGWRD25, UCFGWRD24, UCFGWRD23, UCFGWRD22, UCFGWRD21, UCFGWRD20, UCFGWRD19, UCFGWRD18, UCFGWRD17, UCFGWRD16, UCFGWRD15, UCFGWRD14, UCFGWRD13, UCFGWRD12, UCFGWRD11, UCFGWRD10, UCFGWRD9, UCFGWRD8, UCFGWRD7, UCFGWRD6, UCFGWRD5, UCFGWRD4, UCFGWRD3, UCFGWRD2, UCFGWRD1, UCFGWRD0, UCFGWRDN, USERAUPD, USERTRS3, USERTRS2, USERTRS1, USERTRS0, LMMICLK, LMMIOFFSET16, LMMIOFFSET15, LMMIOFFSET14, LMMIOFFSET13, LMMIOFFSET12, LMMIOFFSET11, LMMIOFFSET10, LMMIOFFSET9, LMMIOFFSET8, LMMIOFFSET7, LMMIOFFSET6, LMMIOFFSET5, LMMIOFFSET4, LMMIOFFSET3, LMMIOFFSET2, LMMIRDATA31, LMMIRDATA30, LMMIRDATA29, LMMIRDATA28, LMMIRDATA27, LMMIRDATA26, LMMIRDATA25, LMMIRDATA24, LMMIRDATA23, LMMIRDATA22, LMMIRDATA21, LMMIRDATA20, LMMIRDATA19, LMMIRDATA18, LMMIRDATA17, LMMIRDATA16, LMMIRDATA15, LMMIRDATA14, LMMIRDATA13, LMMIRDATA12, LMMIRDATA11, LMMIRDATA10, LMMIRDATA9, LMMIRDATA8, LMMIRDATA7, LMMIRDATA6, LMMIRDATA5, LMMIRDATA4, LMMIRDATA3, LMMIRDATA2, LMMIRDATA1, LMMIRDATA0, LMMIRDATAVALID, LMMIREADY, LMMIREQUEST, LMMIRESETN, LMMIWDATA31, LMMIWDATA30, LMMIWDATA29, LMMIWDATA28, LMMIWDATA27, LMMIWDATA26, LMMIWDATA25, LMMIWDATA24, LMMIWDATA23, LMMIWDATA22, LMMIWDATA21, LMMIWDATA20, LMMIWDATA19, LMMIWDATA18, LMMIWDATA17, LMMIWDATA16, LMMIWDATA15, LMMIWDATA14, LMMIWDATA13, LMMIWDATA12, LMMIWDATA11, LMMIWDATA10, LMMIWDATA9, LMMIWDATA8, LMMIWDATA7, LMMIWDATA6, LMMIWDATA5, LMMIWDATA4, LMMIWDATA3, LMMIWDATA2, LMMIWDATA1, LMMIWDATA0, LMMIWRRDN, VRXCMDD12, VRXCMDD11, VRXCMDD10, VRXCMDD9, VRXCMDD8, VRXCMDD7, VRXCMDD6, VRXCMDD5, VRXCMDD4, VRXCMDD3, VRXCMDD2, VRXCMDD1, VRXCMDD0, VRXCINIT, VRXCNH11, VRXCNH10, VRXCNH9, VRXCNH8, VRXCNH7, VRXCNH6, VRXCNH5, VRXCNH4, VRXCNH3, VRXCNH2, VRXCNH1, VRXCNH0, VRXCNINF, VRXCRRE, VRXD31, VRXD30, VRXD29, VRXD28, VRXD27, VRXD26, VRXD25, VRXD24, VRXD23, VRXD22, VRXD21, VRXD20, VRXD19, VRXD18, VRXD17, VRXD16, VRXD15, VRXD14, VRXD13, VRXD12, VRXD11, VRXD10, VRXD9, VRXD8, VRXD7, VRXD6, VRXD5, VRXD4, VRXD3, VRXD2, VRXD1, VRXD0, VRXDP3, VRXDP2, VRXDP1, VRXDP0, VRXEOP, VRXERR, VRXF1, VRXF0, VRXRDY, VRXSEL1, VRXSEL0, VRXSOP, VRXVD, VXCDINIT, VXCDNH11, VXCDNH10, VXCDNH9, VXCDNH8, VXCDNH7, VXCDNH6, VXCDNH5, VXCDNH4, VXCDNH3, VXCDNH2, VXCDNH1, VXCDNH0, VTXCRRE, VXD31, VXD30, VXD29, VXD28, VXD27, VXD26, VXD25, VXD24, VXD23, VXD22, VXD21, VXD20, VXD19, VXD18, VXD17, VXD16, VXD15, VXD14, VXD13, VXD12, VXD11, VXD10, VXD9, VXD8, VXD7, VXD6, VXD5, VXD4, VXD3, VXD2, VXD1, VXD0, VXDP3, VXDP2, VXDP1, VXDP0, VXEOP, VXEOPN, VXRDY, VXSOP, VXVD, TESTOUT7, TESTOUT6, TESTOUT5, TESTOUT4, TESTOUT3, TESTOUT2, TESTOUT1, TESTOUT0, REFCLKNA, S0REFCKN, S0REFCKP, S0REFRET, S0REXT, S0RXN, S0RXP, S0TXN, S0TXP, CLKREQI, CLKREQO, CLKREQOE, SCANCLK, SCANRST, OPCGLDCK, ALTCLKIN); //synthesis syn_black_box black_box_pad_pin="S0REFCKN,S0REFCKP,S0REFRET,S0REXT,S0RXN,S0RXP,S0TXN,S0TXP" syn_lib_cell=1

	input ACTACMD;
	input ACTDR11;
	input ACTEN;
	input ACTHIGHZ;
	input ACTMD;
	output ACJNOUT;
	output ACJPOUT;
	input AUXCK;
	input CKUSRI;
	output CKUSRO;
	input ECKIN;
	input ECKIND2;
	output ECKINDO;
	input ERSTN;
	input ERSTND2;
	input ERXCKD2;
	output ERXCKDO;
	input ERXRSND2;
	input ETXCKD2;
	output ETXCKDO;
	input ETXRSND2;
	output FLR3;
	output FLR2;
	output FLR1;
	output FLR0;
	input FLRACK3;
	input FLRACK2;
	input FLRACK1;
	input FLRACK0;
	input MINTLEG3;
	input MINTLEG2;
	input MINTLEG1;
	input MINTLEG0;
	output MINTO;
	input PERSTN;
	output PMCTRL4;
	output PMCTRL3;
	output PMCTRL2;
	output PMCTRL1;
	output PMCTRL0;
	output PMCTRLEN;
	input PMDPAST4;
	input PMDPAST3;
	input PMDPAST2;
	input PMDPAST1;
	input PMDPAST0;
	input PRMSGSD;
	input PRNOSNP12;
	input PRNOSNP11;
	input PRNOSNP10;
	input PRNOSNP9;
	input PRNOSNP8;
	input PRNOSNP7;
	input PRNOSNP6;
	input PRNOSNP5;
	input PRNOSNP4;
	input PRNOSNP3;
	input PRNOSNP2;
	input PRNOSNP1;
	input PRNOSNP0;
	input PRNSNPRE;
	input PRSNOOP12;
	input PRSNOOP11;
	input PRSNOOP10;
	input PRSNOOP9;
	input PRSNOOP8;
	input PRSNOOP7;
	input PRSNOOP6;
	input PRSNOOP5;
	input PRSNOOP4;
	input PRSNOOP3;
	input PRSNOOP2;
	input PRSNOOP1;
	input PRSNOOP0;
	input PRSNPRE;
	input PPBDREG31;
	input PPBDREG30;
	input PPBDREG29;
	input PPBDREG28;
	input PPBDREG27;
	input PPBDREG26;
	input PPBDREG25;
	input PPBDREG24;
	input PPBDREG23;
	input PPBDREG22;
	input PPBDREG21;
	input PPBDREG20;
	input PPBDREG19;
	input PPBDREG18;
	input PPBDREG17;
	input PPBDREG16;
	input PPBDREG15;
	input PPBDREG14;
	input PPBDREG13;
	input PPBDREG12;
	input PPBDREG11;
	input PPBDREG10;
	input PPBDREG9;
	input PPBDREG8;
	input PPBDREG7;
	input PPBDREG6;
	input PPBDREG5;
	input PPBDREG4;
	input PPBDREG3;
	input PPBDREG2;
	input PPBDREG1;
	input PPBDREG0;
	output PPBDSEL7;
	output PPBDSEL6;
	output PPBDSEL5;
	output PPBDSEL4;
	output PPBDSEL3;
	output PPBDSEL2;
	output PPBDSEL1;
	output PPBDSEL0;
	input REXTCK;
	input REXTRST;
	input RSTUSRN;
	output UDLLKUP;
	input ULTSDIS;
	output UPLLKUP;
	output UTLLKUP;
	input UCFGADDR11;
	input UCFGADDR10;
	input UCFGADDR9;
	input UCFGADDR8;
	input UCFGADDR7;
	input UCFGADDR6;
	input UCFGADDR5;
	input UCFGADDR4;
	input UCFGADDR3;
	input UCFGADDR2;
	input UCFGF2;
	input UCFGF1;
	input UCFGF0;
	output UCFGRDD31;
	output UCFGRDD30;
	output UCFGRDD29;
	output UCFGRDD28;
	output UCFGRDD27;
	output UCFGRDD26;
	output UCFGRDD25;
	output UCFGRDD24;
	output UCFGRDD23;
	output UCFGRDD22;
	output UCFGRDD21;
	output UCFGRDD20;
	output UCFGRDD19;
	output UCFGRDD18;
	output UCFGRDD17;
	output UCFGRDD16;
	output UCFGRDD15;
	output UCFGRDD14;
	output UCFGRDD13;
	output UCFGRDD12;
	output UCFGRDD11;
	output UCFGRDD10;
	output UCFGRDD9;
	output UCFGRDD8;
	output UCFGRDD7;
	output UCFGRDD6;
	output UCFGRDD5;
	output UCFGRDD4;
	output UCFGRDD3;
	output UCFGRDD2;
	output UCFGRDD1;
	output UCFGRDD0;
	output UCFGRDE;
	output UCFGRDY;
	input UCFGSERD;
	input UCFGVD;
	input UCFGWRBE3;
	input UCFGWRBE2;
	input UCFGWRBE1;
	input UCFGWRBE0;
	input UCFGWRD31;
	input UCFGWRD30;
	input UCFGWRD29;
	input UCFGWRD28;
	input UCFGWRD27;
	input UCFGWRD26;
	input UCFGWRD25;
	input UCFGWRD24;
	input UCFGWRD23;
	input UCFGWRD22;
	input UCFGWRD21;
	input UCFGWRD20;
	input UCFGWRD19;
	input UCFGWRD18;
	input UCFGWRD17;
	input UCFGWRD16;
	input UCFGWRD15;
	input UCFGWRD14;
	input UCFGWRD13;
	input UCFGWRD12;
	input UCFGWRD11;
	input UCFGWRD10;
	input UCFGWRD9;
	input UCFGWRD8;
	input UCFGWRD7;
	input UCFGWRD6;
	input UCFGWRD5;
	input UCFGWRD4;
	input UCFGWRD3;
	input UCFGWRD2;
	input UCFGWRD1;
	input UCFGWRD0;
	input UCFGWRDN;
	input USERAUPD;
	input USERTRS3;
	input USERTRS2;
	input USERTRS1;
	input USERTRS0;
	input LMMICLK;
	input LMMIOFFSET16;
	input LMMIOFFSET15;
	input LMMIOFFSET14;
	input LMMIOFFSET13;
	input LMMIOFFSET12;
	input LMMIOFFSET11;
	input LMMIOFFSET10;
	input LMMIOFFSET9;
	input LMMIOFFSET8;
	input LMMIOFFSET7;
	input LMMIOFFSET6;
	input LMMIOFFSET5;
	input LMMIOFFSET4;
	input LMMIOFFSET3;
	input LMMIOFFSET2;
	output LMMIRDATA31;
	output LMMIRDATA30;
	output LMMIRDATA29;
	output LMMIRDATA28;
	output LMMIRDATA27;
	output LMMIRDATA26;
	output LMMIRDATA25;
	output LMMIRDATA24;
	output LMMIRDATA23;
	output LMMIRDATA22;
	output LMMIRDATA21;
	output LMMIRDATA20;
	output LMMIRDATA19;
	output LMMIRDATA18;
	output LMMIRDATA17;
	output LMMIRDATA16;
	output LMMIRDATA15;
	output LMMIRDATA14;
	output LMMIRDATA13;
	output LMMIRDATA12;
	output LMMIRDATA11;
	output LMMIRDATA10;
	output LMMIRDATA9;
	output LMMIRDATA8;
	output LMMIRDATA7;
	output LMMIRDATA6;
	output LMMIRDATA5;
	output LMMIRDATA4;
	output LMMIRDATA3;
	output LMMIRDATA2;
	output LMMIRDATA1;
	output LMMIRDATA0;
	output LMMIRDATAVALID;
	output LMMIREADY;
	input LMMIREQUEST;
	input LMMIRESETN;
	input LMMIWDATA31;
	input LMMIWDATA30;
	input LMMIWDATA29;
	input LMMIWDATA28;
	input LMMIWDATA27;
	input LMMIWDATA26;
	input LMMIWDATA25;
	input LMMIWDATA24;
	input LMMIWDATA23;
	input LMMIWDATA22;
	input LMMIWDATA21;
	input LMMIWDATA20;
	input LMMIWDATA19;
	input LMMIWDATA18;
	input LMMIWDATA17;
	input LMMIWDATA16;
	input LMMIWDATA15;
	input LMMIWDATA14;
	input LMMIWDATA13;
	input LMMIWDATA12;
	input LMMIWDATA11;
	input LMMIWDATA10;
	input LMMIWDATA9;
	input LMMIWDATA8;
	input LMMIWDATA7;
	input LMMIWDATA6;
	input LMMIWDATA5;
	input LMMIWDATA4;
	input LMMIWDATA3;
	input LMMIWDATA2;
	input LMMIWDATA1;
	input LMMIWDATA0;
	input LMMIWRRDN;
	output VRXCMDD12;
	output VRXCMDD11;
	output VRXCMDD10;
	output VRXCMDD9;
	output VRXCMDD8;
	output VRXCMDD7;
	output VRXCMDD6;
	output VRXCMDD5;
	output VRXCMDD4;
	output VRXCMDD3;
	output VRXCMDD2;
	output VRXCMDD1;
	output VRXCMDD0;
	input VRXCINIT;
	input VRXCNH11;
	input VRXCNH10;
	input VRXCNH9;
	input VRXCNH8;
	input VRXCNH7;
	input VRXCNH6;
	input VRXCNH5;
	input VRXCNH4;
	input VRXCNH3;
	input VRXCNH2;
	input VRXCNH1;
	input VRXCNH0;
	input VRXCNINF;
	input VRXCRRE;
	output VRXD31;
	output VRXD30;
	output VRXD29;
	output VRXD28;
	output VRXD27;
	output VRXD26;
	output VRXD25;
	output VRXD24;
	output VRXD23;
	output VRXD22;
	output VRXD21;
	output VRXD20;
	output VRXD19;
	output VRXD18;
	output VRXD17;
	output VRXD16;
	output VRXD15;
	output VRXD14;
	output VRXD13;
	output VRXD12;
	output VRXD11;
	output VRXD10;
	output VRXD9;
	output VRXD8;
	output VRXD7;
	output VRXD6;
	output VRXD5;
	output VRXD4;
	output VRXD3;
	output VRXD2;
	output VRXD1;
	output VRXD0;
	output VRXDP3;
	output VRXDP2;
	output VRXDP1;
	output VRXDP0;
	output VRXEOP;
	output VRXERR;
	output VRXF1;
	output VRXF0;
	input VRXRDY;
	output VRXSEL1;
	output VRXSEL0;
	output VRXSOP;
	output VRXVD;
	output VXCDINIT;
	output VXCDNH11;
	output VXCDNH10;
	output VXCDNH9;
	output VXCDNH8;
	output VXCDNH7;
	output VXCDNH6;
	output VXCDNH5;
	output VXCDNH4;
	output VXCDNH3;
	output VXCDNH2;
	output VXCDNH1;
	output VXCDNH0;
	output VTXCRRE;
	input VXD31;
	input VXD30;
	input VXD29;
	input VXD28;
	input VXD27;
	input VXD26;
	input VXD25;
	input VXD24;
	input VXD23;
	input VXD22;
	input VXD21;
	input VXD20;
	input VXD19;
	input VXD18;
	input VXD17;
	input VXD16;
	input VXD15;
	input VXD14;
	input VXD13;
	input VXD12;
	input VXD11;
	input VXD10;
	input VXD9;
	input VXD8;
	input VXD7;
	input VXD6;
	input VXD5;
	input VXD4;
	input VXD3;
	input VXD2;
	input VXD1;
	input VXD0;
	input VXDP3;
	input VXDP2;
	input VXDP1;
	input VXDP0;
	input VXEOP;
	input VXEOPN;
	output VXRDY;
	input VXSOP;
	input VXVD;
	output TESTOUT7;
	output TESTOUT6;
	output TESTOUT5;
	output TESTOUT4;
	output TESTOUT3;
	output TESTOUT2;
	output TESTOUT1;
	output TESTOUT0;
	input REFCLKNA;
	input S0REFCKN;
	input S0REFCKP;
	input S0REFRET;
	input S0REXT;
	input S0RXN;
	input S0RXP;
	output S0TXN;
	output S0TXP;
	input CLKREQI;
	output CLKREQO;
	output CLKREQOE;
	input SCANCLK;
	input SCANRST;
	input OPCGLDCK;
	input ALTCLKIN;

	parameter ENABLE_USER_CFG = "DISABLED";
	parameter PWDN_N = "DISABLED";
	parameter GSR = "ENABLED";
	parameter IDDQ_PCS = "DISABLED";
	parameter PHY_MODE = "0b0000";
	parameter ALT_CLK_SEL_VCC = "PAD";
	parameter L0S_ADJ = "0b00000110000000";
	parameter L0S_EXIT_LATENCY = "MORE_4_US";
	parameter L1_EXIT_LATENCY = "MORE_64_US";
	parameter CALIB_3DB = "ENABLED";
	parameter DB_UPSTREAM = "6DB";
	parameter ERR_REC_ENTRY_SEL = "RCVRY_AFTER";
	parameter A_CHNGD_MAX = "0b100";
	parameter A0_FORCE = "DISABLED";
	parameter A0_FREEZE = "DISABLED";
	parameter A0_INIT = "0b000000";
	parameter A0DIR_VAL = "DISABLED";
	parameter A1_FORCE = "DISABLED";
	parameter A1_FREEZE = "DISABLED";
	parameter A1_INIT = "0b000000";
	parameter A1DIR_VAL = "DISABLED";
	parameter A2_FORCE = "DISABLED";
	parameter A2_FREEZE = "DISABLED";
	parameter A2_INIT = "0b000000";
	parameter A2GAIN_CALIB = "0b100110";
	parameter ACJTAG_REG = "0b00";
	parameter ADDR_LIMIT_PRE_MTHD_CTRL = "0b0100";
	parameter ADDR_LIMIT_TABLE_MTHD_CTRL = "0b00101";
	parameter ADIR_OVR = "DISABLED";
	parameter ADV_CH_CD_SEL = "IMPLEMENT_CH";
	parameter ADV_TARGET_LINK_SPEED_USPORT_A = "DISABLED";
	parameter ADV_TARGET_LINK_SPEED_USPORT_B = "DISABLED";
	parameter ADV_TARGET_LINK_SPEED_USPORT_C = "DISABLED";
	parameter ADV_TARGET_LINK_SPEED_USPORT_D = "DISABLED";
	parameter ADVANCE = "DISABLED";
	parameter ALERT_ENABLE = "0b000";
	parameter ALMOST_EMPTY_10B = "0b001110";
	parameter MID_VALUE_10B = "0b011110";
	parameter ALMOST_EMPTY_20B = "0b001111";
	parameter ALMOST_EMPTY_GEN3 = "0b001100";
	parameter ALMOST_FULL_10B = "0b110000";
	parameter ALMOST_FULL_20B = "0b011000";
	parameter ALMOST_FULL_GEN3 = "0b010110";
	parameter ARRAY_DA = "0b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter ARRAY_MT = "0b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000011100000000000010000000000000001001000000000000011000000000000001010000000000000100";
	parameter ARXCDRICP_RATE0 = "0b011";
	parameter ARXCDRICP_RATE1 = "0b011";
	parameter ARXCDRICP_RATE2 = "0b011";
	parameter ARXDMPWRDWN = "DISABLED";
	parameter ARXDPPWRDN = "DISABLED";
	parameter ARXEOM_PWRDN = "POWERED_DOWN";
	parameter ARXICP_RATE0 = "0b011";
	parameter ARXICP_RATE1 = "0b011";
	parameter ARXICP_RATE2 = "0b011";
	parameter ARXOVR_OUT = "DISABLED";
	parameter ARXRSACTAT = "0b0001";
	parameter ARXRSAPTAT = "0b1000";
	parameter ARXRSVCTL = "0b00000000";
	parameter ARXSEL_OUT = "DISABLED";
	parameter ASPM_L1_1_SUPPORTED = "SUPPORTED";
	parameter ASPM_L1_2_SUPPORTED = "SUPPORTED";
	parameter ASPM_SUPPORT = "L0S_AND_L1_SUPPORTED";
	parameter ATTENTION_BUTTON_PRESENT = "NOT_SUPPORTED";
	parameter ATTENTION_INDICATOR_PRESENT = "NOT_SUPPORTED";
	parameter ATXICP_RATE0 = "0b101";
	parameter ATXICP_RATE1 = "0b101";
	parameter AUTO_SHIFT = "ENABLED";
	parameter AUX_CURRENT = "SELF_POWERED";
	parameter AUXCLK1US_MAX = "0b00001001";
	parameter AUXIDL_MAX = "0b00000100";
	parameter BAR_INDEX_CFG0_A = "0b000";
	parameter BAR_INDEX_CFG0_B = "0b000";
	parameter BAR_INDEX_CFG0_C = "0b000";
	parameter BAR_INDEX_CFG0_D = "0b000";
	parameter BAR_INDEX_CFG1_A = "0b001";
	parameter BAR_INDEX_CFG1_B = "0b001";
	parameter BAR_INDEX_CFG1_C = "0b001";
	parameter BAR_INDEX_CFG1_D = "0b001";
	parameter BAR_INDEX_CFG2_A = "0b010";
	parameter BAR_INDEX_CFG2_B = "0b010";
	parameter BAR_INDEX_CFG2_C = "0b010";
	parameter BAR_INDEX_CFG2_D = "0b010";
	parameter BAR_INDEX_CFG3_A = "0b011";
	parameter BAR_INDEX_CFG3_B = "0b011";
	parameter BAR_INDEX_CFG3_C = "0b011";
	parameter BAR_INDEX_CFG3_D = "0b011";
	parameter BAR_INDEX_CFG4_A = "0b100";
	parameter BAR_INDEX_CFG4_B = "0b100";
	parameter BAR_INDEX_CFG4_C = "0b100";
	parameter BAR_INDEX_CFG4_D = "0b100";
	parameter BAR_INDEX_CFG5_A = "0b101";
	parameter BAR_INDEX_CFG5_B = "0b101";
	parameter BAR_INDEX_CFG5_C = "0b101";
	parameter BAR_INDEX_CFG5_D = "0b101";
	parameter BIR_MSIX_PBA_A = "BAR0";
	parameter BIR_MSIX_PBA_B = "BAR0";
	parameter BIR_MSIX_PBA_C = "BAR0";
	parameter BIR_MSIX_PBA_D = "BAR0";
	parameter BIR_MSIX_TABLE_A = "BAR0";
	parameter BIR_MSIX_TABLE_B = "BAR0";
	parameter BIR_MSIX_TABLE_C = "BAR0";
	parameter BIR_MSIX_TABLE_D = "BAR0";
	parameter BYP_AVG = "USED";
	parameter BYPASS = "PERFORM_RECEIVER_DETECTION";
	parameter BYPASS_ADDR_DEC = "NORMAL";
	parameter CALIB_SETTLE_MAX = "0b001";
	parameter CALIB_STABLE_MAX = "0b11000";
	parameter CAPABILITY_VERSION = "0b0010";
	parameter CDR_ERR = "DISABLED";
	parameter CDR_P1 = "CDR_PLL_RESET";
	parameter CDR_PLL_DELTA = "0P4_PERCENT";
	parameter CDR_REFERENCE = "0b00";
	parameter CDRPLL_CMP_MAX = "0b00010100";
	parameter CDRPLL_CNT_MAX = "0b00000100";
	parameter CDRPLL_PRE_RXEQ_COARSE_TIMER = "0b01010000";
	parameter CDRPLL_PRE_RXEQ_FINE_TIMER = "0b10110100";
	parameter CDRPLL_PST_RXEQ_COARSE_TIMER = "0b01000000";
	parameter CDRPLL_PST_RXEQ_FINE_TIMER = "0b01000010";
	parameter CFG_A_BAR0 = "0b11111111111111110000000000001100";
	parameter CFG_A_BAR1 = "0b11111111111111111111111111111111";
	parameter CFG_A_BAR2 = "0b11111111111111111110000000001100";
	parameter CFG_A_BAR3 = "0b11111111111111111111111111111111";
	parameter CFG_A_BAR4 = "0b11111111111111111110000000001100";
	parameter CFG_A_BAR5 = "0b11111111111111111111111111111111";
	parameter CFG_B_BAR0 = "0b11111111111111110000000000001100";
	parameter CFG_B_BAR1 = "0b11111111111111111111111111111111";
	parameter CFG_B_BAR2 = "0b11111111111111111110000000001100";
	parameter CFG_B_BAR3 = "0b11111111111111111111111111111111";
	parameter CFG_B_BAR4 = "0b11111111111111111110000000001100";
	parameter CFG_B_BAR5 = "0b11111111111111111111111111111111";
	parameter CFG_C_BAR0 = "0b11111111111111110000000000001100";
	parameter CFG_C_BAR1 = "0b11111111111111111111111111111111";
	parameter CFG_C_BAR2 = "0b11111111111111111110000000001100";
	parameter CFG_C_BAR3 = "0b11111111111111111111111111111111";
	parameter CFG_C_BAR4 = "0b11111111111111111110000000001100";
	parameter CFG_C_BAR5 = "0b11111111111111111111111111111111";
	parameter CFG_D_BAR0 = "0b11111111111111110000000000001100";
	parameter CFG_D_BAR1 = "0b11111111111111111111111111111111";
	parameter CFG_D_BAR2 = "0b11111111111111111110000000001100";
	parameter CFG_D_BAR3 = "0b11111111111111111111111111111111";
	parameter CFG_D_BAR4 = "0b11111111111111111110000000001100";
	parameter CFG_D_BAR5 = "0b11111111111111111111111111111111";
	parameter CFG_EXP_ROM_A = "0b00000000000000000000000000000000";
	parameter CFG_EXP_ROM_B = "0b00000000000000000000000000000000";
	parameter CFG_EXP_ROM_C = "0b00000000000000000000000000000000";
	parameter CFG_EXP_ROM_D = "0b00000000000000000000000000000000";
	parameter CIS_POINTER_CARDBUS_A = "0b00000000000000000000000000000000";
	parameter CIS_POINTER_CARDBUS_B = "0b00000000000000000000000000000000";
	parameter CIS_POINTER_CARDBUS_C = "0b00000000000000000000000000000000";
	parameter CIS_POINTER_CARDBUS_D = "0b00000000000000000000000000000000";
	parameter CLASS_CODE_ID3A = "0b000100011000000000000000";
	parameter CLASS_CODE_ID3B = "0b000100011000000000000000";
	parameter CLASS_CODE_ID3C = "0b000100011000000000000000";
	parameter CLASS_CODE_ID3D = "0b000100011000000000000000";
	parameter CM_RESTORE_TIME = "0b00000000";
	parameter CNT250NS_MAX = "0b001111100";
	parameter COARSE_GAIN = "DISABLED";
	parameter COEF_EN_LPBK_MASTER = "OTHERWISE";
	parameter COEF_EN_LPBK_SLAVE = "OTHERWISE";
	parameter COEF_ENABLE = "DETERMINE_LOCAL_PHY";
	parameter COEF_EQTX_FORCE = "0b000000000000000000";
	parameter COEF_LPBK_MASTER = "0b000000000000000000";
	parameter COEF_LPBK_SLAVE = "0b000000000000000000";
	parameter COEF0_POST = "0b000101";
	parameter COEF0_POST_CURSOR = "0b000000";
	parameter COEF0_PRE = "0b000000";
	parameter COEF0_PRE_CURSOR = "0b000000";
	parameter COEF1_POST = "0b000011";
	parameter COEF1_POST_CURSOR = "0b000000";
	parameter COEF1_PRE = "0b000000";
	parameter COEF1_PRE_CURSOR = "0b000000";
	parameter COEF10_POST = "0b000111";
	parameter COEF10_PRE = "0b000000";
	parameter COEF2_POST = "0b000100";
	parameter COEF2_POST_CURSOR = "0b000000";
	parameter COEF2_PRE = "0b000000";
	parameter COEF2_PRE_CURSOR = "0b000000";
	parameter COEF3_POST = "0b000010";
	parameter COEF3_POST_CURSOR = "0b000000";
	parameter COEF3_PRE = "0b000000";
	parameter COEF3_PRE_CURSOR = "0b000000";
	parameter COEF4_POST = "0b000000";
	parameter COEF4_PRE = "0b000000";
	parameter COEF5_POST = "0b000000";
	parameter COEF5_PRE = "0b000001";
	parameter COEF6_POST = "0b000000";
	parameter COEF6_PRE = "0b000010";
	parameter COEF7_POST = "0b000100";
	parameter COEF7_PRE = "0b000011";
	parameter COEF8_POST = "0b000011";
	parameter COEF8_PRE = "0b000010";
	parameter COEF9_POST = "0b000000";
	parameter COEF9_PRE = "0b000011";
	parameter COMP_128_SUPPORTED = "ENABLED";
	parameter COMP_32_SUPPORTED = "ENABLED";
	parameter COMP_64_SUPPORTED = "ENABLED";
	parameter COMPLETE = "DISABLED";
	parameter CONV_METHOD = "COMPUTE_PCIE_SPEC";
	parameter CORE_BYPASS = "NORMAL";
	parameter CORE_EN = "ENABLED";
	parameter COUNT_ACK_TO_NAK = "0b00000000";
	parameter CPL_TIMEOUT_DISABLE_SUPPORTED = "SUPPORTED";
	parameter CPL_TIMEOUT_RANGES_SUPPORTED = "NOT_SUPPORTED";
	parameter CRS_ENABLE = "DISABLED";
	parameter CSTAT_DATA_SCALE = "UNKNOWN_SCALE";
	parameter CSTAT_DATA_SELECT = "D0_POWER_CONSUMED";
	parameter CTLE_SETTLE = "0b100";
	parameter CTLEBIAS_1 = "0b1000";
	parameter ATXICP_RATE2 = "0b100";
	parameter CTLEBYPASS = "DISABLED";
	parameter CUR_FOM = "NUMBER_OF_CLOCK";
	parameter CUR_FOM_AVG = "0b101";
	parameter CUST_AUTO = "DISABLED";
	parameter CUST_CHK = "SET";
	parameter CUST_SEL = "DISABLED";
	parameter CUST_SKIP = "DISABLED";
	parameter CUST_TYP = "0b000";
	parameter CUSTOM_PATTERN = "0b00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter D1_SUPPORT = "SUPPORTED";
	parameter D2_SUPPORT = "SUPPORTED";
	parameter DATA_INJECT = "0b00000000000000000000000000000000";
	parameter DATA_PM = "0b00000000";
	parameter DEEMPH_5G_3_5DB_6DB_N = "6DB";
	parameter DEEMPH_5G_ENABLE = "DISABLED";
	parameter DEEMPH_LPBK_MASTER = "6P0DB";
	parameter DEEMPH_LPBK_SLAVE = "6P0DB";
	parameter DEVICE_ID_ID1A = "0b1110000000000100";
	parameter DEVICE_ID_ID1B = "0b1110000000000100";
	parameter DEVICE_ID_ID1C = "0b1110000000000100";
	parameter DEVICE_ID_ID1D = "0b1110000000000100";
	parameter DEVICE_PORT_TYPE = "PCIE_ENDPOINT";
	parameter DFE_BIAS = "0b0001";
	parameter DFE_PWDN = "DISABLED";
	parameter DIR_PRE_GAIN = "0b00";
	parameter DIR_PST_GAIN = "0b01";
	parameter DIS_ARI_CAP = "ENABLED";
	parameter DIS_CSR_RST = "DISABLED";
	parameter DIS_INTERRUPT = "ENABLED";
	parameter DIS_INTERRUPT_B = "ENABLED";
	parameter DIS_INTERRUPT_C = "ENABLED";
	parameter DIS_INTERRUPT_D = "ENABLED";
	parameter DIS_MSI_CAP = "ENABLED";
	parameter DIS_MSI_CAP_B = "ENABLED";
	parameter DIS_MSI_CAP_C = "ENABLED";
	parameter DIS_MSI_CAP_D = "ENABLED";
	parameter DIS_MSIX_CAP = "ENABLED";
	parameter DIS_MSIX_CAP_B = "ENABLED";
	parameter DIS_MSIX_CAP_C = "ENABLED";
	parameter DIS_MSIX_CAP_D = "ENABLED";
	parameter DISABLE_FLR_CAPABILITY = "ENABLED";
	parameter DLLP_CRC_ERR_ENABLE = "DISABLED";
	parameter DLLP_CRC_ERR_RATE = "0b000000000000";
	parameter DLLP_INJECT_ENABLE = "DISABLED";
	parameter DOUBLE_TX_DATA_VALID = "ONE_CLK_EVERY_64_CLKS";
	parameter DOWNSTREAM_EQ_SKIP_PHASE_2_3 = "NORMAL_OPERATION";
	parameter DS_DRIVE_CLKREQ = "ENABLED";
	parameter DS_PORT_RX_PRESET_HINT = "0b001";
	parameter DS_PORT_TX_PRESET = "0b0011";
	parameter DS_US_N_PORTTYPE = "UPSTREAM";
	parameter DSI = "NO_DSI_NECESSARY";
	parameter DSP_DIR = "ANALYSIS_OF_DATA_BY_DSP";
	parameter DSPDIR_PRESGN = "0b11110000";
	parameter DSPDIR_PREVAL = "0b00011000";
	parameter DSPDIR_PSTSGN0 = "0b11111111";
	parameter DSPDIR_PSTSGN1 = "0b00000000";
	parameter DSPDIR_PSTVAL0 = "0b00000010";
	parameter DSPDIR_PSTVAL1 = "0b01000000";
	parameter EARLY_RX_EVAL = "RX_SIGNAL_AFTER_TS1";
	parameter ECRC_GEN_CHK_CAPABLE = "SUPPORTED";
	parameter EFF_LPBK = "PASSED";
	parameter EI4 = "EI_IV";
	parameter EM_INTERLOCK_PRESENT = "NOT_SUPPORTED";
	parameter EN = "DISABLED";
	parameter EN_ACK_TO_DIV = "ACK_SPEC";
	parameter EN_ACK_TO_NAK = "DO_NOTHING";
	parameter EN_ACS_VIOLATION = "DISABLED";
	parameter EN_ASPM_L0S = "ENABLED";
	parameter EN_ASPM_L1 = "ENABLED";
	parameter EN_ATOMIC_OP_CAP = "ENABLED";
	parameter EN_ATOMICOP_EGRESS_BLOCKED = "DISABLED";
	parameter EN_ATS_CAP = "ENABLED";
	parameter EN_BDGT_CAP = "DISABLED";
	parameter EN_CAP = "ENABLED";
	parameter EN_CAP_B = "ENABLED";
	parameter EN_CAP_C = "ENABLED";
	parameter EN_CAP_D = "ENABLED";
	parameter EN_COMPLETER_ABORT = "DISABLED";
	parameter EN_COMPLETION_TIMEOUT = "ENABLED";
	parameter EN_CORR_INTERNAL_ERROR = "DISABLED";
	parameter EN_DPA_CAP = "DISABLED";
	parameter EN_DRCT_SCR_OFF = "OTHERWISE";
	parameter EN_DRCT_TO_LPBK = "OTHERWISE";
	parameter EN_EQTX_OVERRIDE = "PIPE_LOCAL_FS_AND_PIPE_LOCAL_LF";
	parameter EN_FORCE_SCR_OFF_FAST = "OTHERWISE";
	parameter EN_L1 = "ENABLED";
	parameter EN_L1PMSS_CAP = "ENABLED";
	parameter EN_L2 = "ENABLED";
	parameter EN_LPBK_ERR_RST = "MASTER_LPBK_INCREMENT";
	parameter EN_LTR_CAP = "ENABLED";
	parameter EN_MC_BLOCKED_TLP = "DISABLED";
	parameter EN_NWL_VSEC_CAP = "ENABLED";
	parameter EN_PORT_DIS = "DISABLED";
	parameter EN_PORT_INTLEG = "ENABLED";
	parameter EN_RBAR_CAP_A = "ENABLED";
	parameter EN_RBAR_CAP_B = "ENABLED";
	parameter EN_RBAR_CAP_C = "ENABLED";
	parameter EN_RBAR_CAP_D = "ENABLED";
	parameter EN_RECEIVER_OVERFLOW = "DISABLED";
	parameter EN_SELF_XLINK = "OTHERWISE";
	parameter EN_SURPRISE_DOWN_ERROR = "DISABLED";
	parameter EN_TLP_PREFIX_BLOCKED = "DISABLED";
	parameter EN_UCORR_INTERNAL_ERROR = "DISABLED";
	parameter EN_USER_WRITE = "READ_WRITE_ACCESS";
	parameter END_END_PREFIXES_SUPPORTED = "NOT_SUPPORTED";
	parameter END_ON_HOLD = "YES_EXIT_ON_HOLD";
	parameter ENDCALIB_MAX = "0b10000100";
	parameter ENDPOINT_L0S_ACCEPTABLE_LATENCY = "MAX_64_NS";
	parameter ENDPOINT_L1_ACCEPTABLE_LATENCY = "MAX_1_US";
	parameter ENTRY_TIME_ASPM_L0S = "0b0000000000000000";
	parameter ENTRY_TIME_ASPM_L1 = "0b0000000000000000";
	parameter EOM_TIME = "0b0000000000000000";
	parameter EOM0DIR = "SELECT_DIR_1";
	parameter EOM1DIR = "SELECT_DIR_0";
	parameter EOMCTRL0_LOW = "DISABLED";
	parameter EOMDIVDIS = "DISABLED";
	parameter EOMMODE = "0b00";
	parameter EOMRDSEL = "DISABLED";
	parameter EOMSTART = "DISABLED";
	parameter EOMX = "0b000000";
	parameter EOMX_UPDATE_CNT_VALUE = "0b0011111";
	parameter EOMY = "0b00000000";
	parameter ERRCNT_DEC = "0b00100000";
	parameter ERRCNT_THR = "0b1000";
	parameter ES_PWDN = "DISABLED";
	parameter EVAL_RST = "DISABLED";
	parameter EXCLUDE_L0 = "INCLUDE";
	parameter EXCLUDE_CFG_COMPLETE = "INCLUDE";
	parameter EXCLUDE_CFG_IDLE = "INCLUDE";
	parameter EXCLUDE_LOOPBACK_MASTER = "INCLUDE";
	parameter EXCLUDE_REC_IDLE = "INCLUDE";
	parameter EXCLUDE_REC_RCVR_CFG = "INCLUDE";
	parameter EXIT_DIRECT_TO_DETECT = "DO_NOT_EXIT_TO_DETECT";
	parameter EXT_CONTROL = "DISABLED";
	parameter EXTENDED_TAG_FIELD_EN_DEFAULT = "EIGHT_BIT";
	parameter EXTENDED_TAG_FIELD_SUPPORTED = "EIGHT_BIT";
	parameter F_ARXCTLEDIR = "IGNORED";
	parameter F_ARXCTLENULL = "0b0000";
	parameter F_ARXDMDIR = "DISABLED";
	parameter F_ARXDMNULL = "0b00000";
	parameter F_ARXEOMDIR = "IGNORED";
	parameter F_ARXEOMNULL = "0b00000";
	parameter F_ARXESDIR = "IGNORED";
	parameter F_ARXESNULL = "0b00000";
	parameter F_ARXTDIR = "IGNORED";
	parameter F_ARXTNULL = "0b00000";
	parameter F_ASCHCAL = "IGNORED";
	parameter F_ASCHDIR = "IGNORED";
	parameter F_ASCHNULL = "0b0000";
	parameter FAIL_LIMIT_ERR = "RXEQ_NOT_FAIL";
	parameter FAST = "L0";
	parameter FC_UPDATE_TIMER_DISABLE = "ENABLED";
	parameter FC_UPDATE_TIMER_DIV = "PCIE_REC_VALUES";
	parameter FILTER = "0b1001";
	parameter FINE_GAIN = "DISABLED";
	parameter FOM_COMPARE = "0b00000000";
	parameter FOM_HIRES = "DISABLED";
	parameter FOM_ITERCNT = "0b101";
	parameter FOM_THR = "0b0100";
	parameter FORCE_ATXDRA = "0b000000000000000000000";
	parameter FORCE_ATXDRP = "0b000000000000000000000";
	parameter FORCE_ATXDRR = "0b000000000000000000000";
	parameter FORCE_ATXDRT = "0b000000000000000000000";
	parameter FORCE_DIR_RSLT = "0b000000";
	parameter FORCE_FOM_RSLT = "0b00000000";
	parameter FORCE_IDLE = "DISABLED";
	parameter FORCE_RX_DETECT = "DISABLED";
	parameter FORCE_SIGNAL = "DISABLED";
	parameter FREQ_LOCK = "DISABLED";
	parameter FS = "0b110000";
	parameter GAIN_TIMER1 = "0b0101";
	parameter GEN12_ENA_POST_A0 = "DISABLED";
	parameter GEN12_ENA_POST_A1A2 = "DISABLED";
	parameter GEN12_ENA_PREA0 = "DISABLED";
	parameter GEN3_ENA_POST_A0 = "ENABLED";
	parameter GEN3_ENA_POST_A1A2 = "ENABLED";
	parameter GEN3_ENA_PREA0 = "ENABLED";
	parameter GLOBAL_INVAL_SUPPORT = "ENABLED";
	parameter HINT = "0b000";
	parameter HINT0_3DB = "ENABLED";
	parameter HINT0_A0GAIN = "0b111";
	parameter HINT0_A2GAIN = "0b111";
	parameter HINT1_3DB = "ENABLED";
	parameter HINT1_A0GAIN = "0b011";
	parameter HINT1_A2GAIN = "0b101";
	parameter HINT2_3DB = "ENABLED";
	parameter HINT2_A0GAIN = "0b011";
	parameter HINT2_A2GAIN = "0b111";
	parameter HINT3_3DB = "ENABLED";
	parameter HINT3_A0GAIN = "0b000";
	parameter HINT3_A2GAIN = "0b111";
	parameter HINT4_3DB = "DISABLED";
	parameter HINT4_A0GAIN = "0b111";
	parameter HINT4_A2GAIN = "0b111";
	parameter HINT5_3DB = "DISABLED";
	parameter HINT5_A0GAIN = "0b011";
	parameter HINT5_A2GAIN = "0b101";
	parameter HINT6_3DB = "DISABLED";
	parameter HINT6_A0GAIN = "0b011";
	parameter HINT6_A2GAIN = "0b111";
	parameter HINT7_3DB = "DISABLED";
	parameter HINT7_A0GAIN = "0b000";
	parameter HINT7_A2GAIN = "0b111";
	parameter HINT7_OVR = "DISABLED";
	parameter HLD_RST = "WRITE_1";
	parameter HOT_PLUG_CAPABLE = "NOT_SUPPORTED";
	parameter HOT_PLUG_SURPRISE = "NOT_POSSIBLE";
	parameter ID_DS_PORT = "0b0000000000000000";
	parameter ID_NWL_VSEC_CAP = "0b0000000000000001";
	parameter IGNORE_ECRC = "DISABLED";
	parameter IGNORE_POISON = "ENABLED";
	parameter INDICATOR = "0b00000000000000000000000000000000";
	parameter INHIBIT = "PERFORM_RECEIVER_DETECTION";
	parameter INJECT_DATA_ERROR_0 = "DISABLED";
	parameter INJECT_DATA_ERROR_1 = "DISABLED";
	parameter INJECT_DATA_ERROR_2 = "DISABLED";
	parameter INJECT_DATA_ERROR_3 = "DISABLED";
	parameter INJECT_DATA_ERROR_EN = "DISABLED";
	parameter INJECT_ERR_LANE_SELECT_0 = "DISABLED";
	parameter INJECT_ERR_LANE_SELECT_1 = "DISABLED";
	parameter INJECT_ERR_LANE_SELECT_2 = "DISABLED";
	parameter INJECT_ERR_LANE_SELECT_3 = "DISABLED";
	parameter INJECT_RX_1BIT_DATA_ERR = "DISABLED";
	parameter INJECT_RX_2BIT_DATA_ERR = "DISABLED";
	parameter INJECT_RX_SKP_ERR = "DISABLED";
	parameter INJECT_RX_VALID_ERR = "DISABLED";
	parameter INT_CLR = "DISABLED";
	parameter INT_EN = "DISABLED";
	parameter INTERRUPT_MESSAGE_NUMBER = "0b00000";
	parameter INVAL_Q_DEPTH = "0b00000";
	parameter ITERATION_MAX = "0b000000";
	parameter L1_ENTER_PLL_RESET_TIME = "0b100";
	parameter L1_EXIT_PLL_LOCK_TIME = "0b01110";
	parameter L1PM_SUPPORTED = "SUPPORTED";
	parameter L2_D3HOT_ENABLE = "DISABLED";
	parameter LANE_SELECT = "0b0000";
	parameter LF = "0b001000";
	parameter LF_PHY = "0b001010";
	parameter LINK_LANE = "ENABLED";
	parameter LPBK_EN = "DISABLED";
	parameter LW_START_UPDN_ACK_EN = "DISABLED";
	parameter LW_START_UPDN_COUNT = "0b000011111010";
	parameter LW_START_UPDN_EIE_EN = "DISABLED";
	parameter LW_START_UPDN_EN_DIR_DS = "DO_NOT_ASSERT";
	parameter LW_START_UPDN_END_DELAY = "0b1001";
	parameter LW_START_UPDN_RATE_EN_16G = "DISABLED";
	parameter LW_START_UPDN_RATE_EN_2P5G = "ENABLED";
	parameter LW_START_UPDN_RATE_EN_5G = "ENABLED";
	parameter LW_START_UPDN_RATE_EN_8G = "ENABLED";
	parameter LW_START_UPDN_START_DELAY = "0b1000";
	parameter LW_START_UPDN_TIMER_EN = "DISABLED";
	parameter MARGIN_ENABLE = "PCIE_SPEC";
	parameter MARGIN_VALUE = "0b000";
	parameter MASK_0 = "SKIP_RCVR_DETECTION";
	parameter MASK_1 = "SKIP_RCVR_DETECTION";
	parameter MASK_2 = "SKIP_RCVR_DETECTION";
	parameter MASK_3 = "SKIP_RCVR_DETECTION";
	parameter MAX_LINK_WIDTH = "1_LANE";
	parameter MAX_SPEED = "8G";
	parameter MAX_VAR = "0b00100";
	parameter MERGE_LMMI_RDATA = "DISABLED";
	parameter METHOD_FMERIT_CTRL = "STEP_PCIE_TX_PRESETS";
	parameter METHOD_TX_CRED_CLEANUP = "HEADER";
	parameter MGMT_INTLEG = "0b0000";
	parameter MGMT_LTSSM_DIS = "DISABLED";
	parameter MID_VALUE_20B = "0b010100";
	parameter MID_VALUE_GEN3 = "0b001110";
	parameter MIN_SPEED = "2P5G";
	parameter MIN_TIME = "0_MS";
	parameter MIN_TIME_CFG = "4US";
	parameter MIX_DIR = "DISABLED";
	parameter MODE_BFF = "RESTART";
	parameter MRL_SENSOR_PRESENT = "NOT_SUPPORTED";
	parameter MULT_ENABLE = "RECOMMENDED_VALUES";
	parameter MULT_MESSAGE_CAPABLE_MSICAP_A = "EIGHT";
	parameter MULT_MESSAGE_CAPABLE_MSICAP_B = "EIGHT";
	parameter MULT_MESSAGE_CAPABLE_MSICAP_C = "EIGHT";
	parameter MULT_MESSAGE_CAPABLE_MSICAP_D = "EIGHT";
	parameter NFTS = "0b11111111";
	parameter NO_COMMAND_COMPLETED_SUPPORT = "SW_NOTIF_PROVIDED";
	parameter NO_FCMP = "DISABLED";
	parameter NO_REMOTE_CHANGE = "DISABLED";
	parameter NO_TX_IDLE_DELAY = "DATA_VALID_GAP";
	parameter NUM_LANES = "1_LANE";
	parameter NUMBER_DSLINK = "0b00000";
	parameter NUMHI_A = "0b00000000000000000000000000000000";
	parameter NUMHI_B = "0b00000000000000000000000000000000";
	parameter NUMHI_C = "0b00000000000000000000000000000000";
	parameter NUMHI_D = "0b00000000000000000000000000000000";
	parameter NUMHOLD = "SINGLE_HOLD_RESPONSE";
	parameter NUMLO_A = "0b00000000000000000000000000000000";
	parameter NUMLO_B = "0b00000000000000000000000000000000";
	parameter NUMLO_C = "0b00000000000000000000000000000000";
	parameter NUMLO_D = "0b00000000000000000000000000000000";
	parameter OBFF_SUPPORTED = "NOT_SUPPORTED";
	parameter OFFSET_MSIX_PBA_A = "0b00000000000000000111000000000";
	parameter OFFSET_MSIX_PBA_B = "0b00000000000000000111000000000";
	parameter OFFSET_MSIX_PBA_C = "0b00000000000000000111000000000";
	parameter OFFSET_MSIX_PBA_D = "0b00000000000000000111000000000";
	parameter OFFSET_MSIX_TABLE_A = "0b00000000000000000110000000000";
	parameter OFFSET_MSIX_TABLE_B = "0b00000000000000000110000000000";
	parameter OFFSET_MSIX_TABLE_C = "0b00000000000000000110000000000";
	parameter OFFSET_MSIX_TABLE_D = "0b00000000000000000110000000000";
	parameter OVER_CTLE = "DISABLED";
	parameter OVER_RX = "DISABLED";
	parameter OVER_RXDM = "DISABLED";
	parameter OVER_RXDP = "DISABLED";
	parameter OVER_RXES = "DISABLED";
	parameter OVER_RXT = "DISABLED";
	parameter OVER_SCH = "DISABLED";
	parameter OVER_TX = "DISABLED";
	parameter OVERRIDE = "DISABLED";
	parameter OVR_CDR = "DISABLED";
	parameter OVR_DIR = "DISABLED";
	parameter OVR_FOM = "DISABLED";
	parameter OVR_GAIN3DB = "ENABLED";
	parameter OVR_HINT3DB = "ENABLED";
	parameter P_CLK_PERIOD = "0b0000111110100000";
	parameter PAR_LPBK = "DISABLED";
	parameter PAS = "10X";
	parameter PATTERN_0 = "UNSCRAMBLED";
	parameter PATTERN_1 = "UNSCRAMBLED";
	parameter PATTERN_2 = "UNSCRAMBLED";
	parameter PCIPM_L1_1_SUPPORTED = "SUPPORTED";
	parameter PCIPM_L1_2_SUPPORTED = "SUPPORTED";
	parameter PERIOD_SRIS_128B130B = "0b000000";
	parameter PERIOD_SRIS_8B10B = "0b00000000";
	parameter PERIOD_SRNS_128B130B = "0b00000000";
	parameter PERIOD_SRNS_8B10B = "0b00000000";
	parameter PHANTOM_FUNCTIONS_SUPPORTED = "NO_FUNCTION_BITS";
	parameter PHYSICAL_SLOT_NUMBER = "0b0000000000001";
	parameter PIN_INTERRUPT_A = "INTA";
	parameter PIN_INTERRUPT_B = "INTA";
	parameter PIN_INTERRUPT_C = "INTA";
	parameter PIN_INTERRUPT_D = "INTA";
	parameter PIPE_TX_SWING = "FULL_SWING";
	parameter PLESIO_LPBK = "DISABLED";
	parameter PM_REDUCE_TIMEOUTS = "DISABLED";
	parameter PMA_DRIVEN_MODE = "PCS_DRIVEN";
	parameter PMCSR_B2_B3_SUPPORT = "DISABLED";
	parameter PMCSR_BUS_P_C_EN = "DISABLED";
	parameter PME_CLOCK = "DISABLED";
	parameter PME_SUPPORT = "0b11111";
	parameter PMFF_ALL = "DISABLED";
	parameter PORT_CM_RESTORE_TIME = "0b00000000";
	parameter PORT_NUMBER = "0b00000000";
	parameter PORT_TPOWER_ON_SCALE = "2_US";
	parameter PORT_TPOWER_ON_VALUE = "0b00000";
	parameter POST = "0b000000";
	parameter POST_A0COEF = "0b001";
	parameter POST_A1COEF = "0b001";
	parameter POST_A2COEF = "0b001";
	parameter POST_CURSOR_LIMIT = "0b100000";
	parameter POST_CURSOR_STEP_SIZE = "0b001000";
	parameter POST_ITERCNT = "0b100";
	parameter POST_STEP = "STEP_SIZE_4";
	parameter POWER_CONTROLLER_PRESENT = "NOT_SUPPORTED";
	parameter POWER_INDICATOR_PRESENT = "NOT_SUPPORTED";
	parameter POWER_REQUIRED = "AUX_POWER_NOT_REQUIRED";
	parameter PRBS_CHK = "DISABLED";
	parameter PRBS_GEN = "DISABLED";
	parameter PRBS_TYP = "PRBS7";
	parameter PRE = "0b000000";
	parameter PRE_A0COEF = "0b101";
	parameter PRE_A1COEF = "0b101";
	parameter PRE_A2COEF = "0b101";
	parameter PRE_CURSOR_LIMIT = "0b010000";
	parameter PRE_CURSOR_STEP_SIZE = "0b000100";
	parameter PRE_FOM = "ENABLED";
	parameter PRE_FOM_AVG = "0b100";
	parameter PRE_ITERCNT = "0b100";
	parameter PRE_RXEQ_TIMER = "0b00010100";
	parameter PRE_STEP = "STEP_SIZE_2";
	parameter PRESET_COUNT_INI = "0b0000";
	parameter PRESET_EN_LPBK_MASTER = "OTHERWISE";
	parameter PRESET_EN_LPBK_SLAVE = "OTHERWISE";
	parameter PRESET_ENABLE = "NORMAL_OP";
	parameter PRESET_EQTX_FORCE = "0b0000";
	parameter PRESET_LPBK_MASTER = "0b0000";
	parameter PRESET_LPBK_SLAVE_0 = "OTHERWISE";
	parameter PRESET_LPBK_SLAVE_1 = "OTHERWISE";
	parameter PRESET_LPBK_SLAVE_2 = "OTHERWISE";
	parameter PRESET_LPBK_SLAVE_3 = "OTHERWISE";
	parameter PRESET_REJECT = "0b00000000000";
	parameter PRESET0_POSTCURSOR = "0b1000";
	parameter PRESET0_PRECURSOR = "0b0000";
	parameter PRESET1_POSTCURSOR = "0b0101";
	parameter PRESET1_PRECURSOR = "0b0000";
	parameter PRESET10_POSTCURSOR = "0b1010";
	parameter PRESET10_PRECURSOR = "0b0000";
	parameter PRESET2_POSTCURSOR = "0b0110";
	parameter PRESET2_PRECURSOR = "0b0000";
	parameter PRESET3_POSTCURSOR = "0b0100";
	parameter PRESET3_PRECURSOR = "0b0000";
	parameter PRESET4_POSTCURSOR = "0b0000";
	parameter PRESET4_PRECURSOR = "0b0000";
	parameter PRESET5_POSTCURSOR = "0b0000";
	parameter PRESET5_PRECURSOR = "0b0011";
	parameter PRESET6_POSTCURSOR = "0b0000";
	parameter PRESET6_PRECURSOR = "0b0100";
	parameter PRESET7_POSTCURSOR = "0b0110";
	parameter PRESET7_PRECURSOR = "0b0011";
	parameter PRESET8_POSTCURSOR = "0b0100";
	parameter PRESET8_PRECURSOR = "0b0100";
	parameter PRESET9_POSTCURSOR = "0b0000";
	parameter PRESET9_PRECURSOR = "0b0101";
	parameter PS_REENTRY_TIME = "0b00000000";
	parameter RATE = "2P5G";
	parameter RATE_ENABLE = "INITIAL_SPEED_CHANGES";
	parameter RCB = "DISABLED";
	parameter REC_SPD_INFER_EQ_PH0123 = "EXCLUDE_TIME_SPENT";
	parameter REC_SPD_INFER_RCVR_CFG = "EXCLUDE_TIME_SPENT";
	parameter REC_SPD_INFER_RCVR_LOCK = "EXCLUDE_TIME_SPENT";
	parameter DIS_FUNC_B = "ENABLED";
	parameter DIS_FUNC_C = "ENABLED";
	parameter DIS_FUNC_D = "ENABLED";
	parameter REDUCE_TIMEOUTS_LTSSMSIM = "DISABLED";
	parameter REDUCE_TIMEOUTS_SIM = "DISABLED";
	parameter REDUCE_TS1 = "DISABLED";
	parameter REENTRY_DISABLE = "ENABLED";
	parameter REENTRY_TIME = "0b00000000000000";
	parameter REQ_FEEDBACK = "0b00000000";
	parameter RESET_EIEOS_INTERVAL_COUNT = "DISABLED";
	parameter REVISION_ID_ID3A = "0b00000100";
	parameter REVISION_ID_ID3B = "0b00000100";
	parameter REVISION_ID_ID3C = "0b00000100";
	parameter REVISION_ID_ID3D = "0b00000100";
	parameter RL1 = "0b0011";
	parameter RL2 = "0b0101";
	parameter RL3 = "0b0011";
	parameter ROUTING_SUPPORTED = "DISABLED";
	parameter RP_COMPLETER_EN = "DISABLED";
	parameter RSTCDR_ERR = "ENABLED";
	parameter RSTCDR_FRQ = "ENABLED";
	parameter RSTCDR_IDL = "DISABLED";
	parameter RX_BYPASS_DECODE_EN = "ENABLED";
	parameter RX_BYPASS_MSG_DEC = "NORMAL_OPERATION";
	parameter RX_CONVERT_UR_TO_CA = "NORMAL_OPERATION";
	parameter RX_D_ALLOC_C = "0b0000000001100000";
	parameter RX_D_ALLOC_N = "0b0000000000000110";
	parameter RX_D_ALLOC_P = "0b0000000001101100";
	parameter RX_DIV_MODE1 = "0b10";
	parameter RX_DIV_MODE0 = "DIV_2";
	parameter RX_DIV_MODE2 = "0b00";
	parameter RX_DL_ACTIVE_DISABLE = "BLOCK_RECEPTION_TLP";
	parameter RX_EARLY_FORWARD_DISABLE = "FWD_RX_DATA_LL";
	parameter RX_ERR_COR = "DISABLED";
	parameter RX_ERR_UCOR = "DISABLED";
	parameter RX_FORCE_RO = "DISABLED";
	parameter RX_H_ALLOC_C = "0b000000100000";
	parameter RX_H_ALLOC_N = "0b000000001000";
	parameter RX_H_ALLOC_P = "0b000000010000";
	parameter RX_HIZ = "IGNORED";
	parameter RX_IMPED_RATIO = "0b10000000";
	parameter RX_INHIBIT_ACK_NAK = "PROCESS_RCVD_ACK";
	parameter RX_INHIBIT_TLP = "PROCESS_RCVD_TLP";
	parameter RX_LCRC_INJECT_EN = "DO_NOT_INJECT_ERROR";
	parameter RX_MALF_INJECT_EN = "DO_NOT_INJECT_ERROR";
	parameter RX_POLINV = "NORMAL";
	parameter RX_PRIORITY = "DISABLED";
	parameter RX_PRIORITY_N_STARVE_THRESH = "0b00010000";
	parameter RX_PRIORITY_P_STARVE_THRESH = "0b00010000";
	parameter RX_PWRDN = "IGNORED";
	parameter RX_TLP_VALID = "DISABLED";
	parameter RXEQ_ALGO = "0b111";
	parameter RXEQ_ENABLE = "0b100";
	parameter RXEQ_EVAL_MAX = "0b11111111";
	parameter RXEQ_MANUAL = "DISABLED";
	parameter RXEQ_STATE = "0b0000";
	parameter RXF_A = "0b0100";
	parameter RXF_B = "0b0100";
	parameter RXF_C = "0b0100";
	parameter RXHF_CLKDN = "ENABLED";
	parameter RXIDLE_MAX = "0b1111";
	parameter RXIDLE_MAX2 = "0b0000010000000000";
	parameter RXIDLE_MSB = "0b11";
	parameter RXM_A = "0b10";
	parameter RXM_B = "0b01";
	parameter RXM_C = "0b00";
	parameter RXN_A = "0b00100";
	parameter RXN_B = "0b01001";
	parameter RXN_C = "0b01111";
	parameter RXOFF_SETTLE_MAX = "0b011";
	parameter RXOFF_STABLE_MAX = "0b10000";
	parameter RXPLLINIT = "DISABLED";
	parameter RXPLLRST = "SET";
	parameter SELECT_DIR_FOM_N = "FME_METHOD";
	parameter SELECTABLE_DEEMPHASIS = "6P0DB";
	parameter SEQ_NUM = "0b000000000000";
	parameter SIGNAL_DETECT_THRESHOLD = "125_MV";
	parameter SIZE_CFG0_A = "0b00000";
	parameter SIZE_CFG0_B = "0b00000";
	parameter SIZE_CFG0_C = "0b00000";
	parameter SIZE_CFG0_D = "0b00000";
	parameter SIZE_CFG1_A = "0b00000";
	parameter SIZE_CFG1_B = "0b00000";
	parameter SIZE_CFG1_C = "0b00000";
	parameter SIZE_CFG1_D = "0b00000";
	parameter SIZE_CFG2_A = "0b00000";
	parameter SIZE_CFG2_B = "0b00000";
	parameter SIZE_CFG2_C = "0b00000";
	parameter SIZE_CFG2_D = "0b00000";
	parameter SIZE_CFG3_A = "0b00000";
	parameter SIZE_CFG3_B = "0b00000";
	parameter SIZE_CFG3_C = "0b00000";
	parameter SIZE_CFG3_D = "0b00000";
	parameter SIZE_CFG4_A = "0b00000";
	parameter SIZE_CFG4_B = "0b00000";
	parameter SIZE_CFG4_C = "0b00000";
	parameter SIZE_CFG4_D = "0b00000";
	parameter SIZE_CFG5_A = "0b00000";
	parameter SIZE_CFG5_B = "0b00000";
	parameter SIZE_CFG5_C = "0b00000";
	parameter SIZE_CFG5_D = "0b00000";
	parameter SKIP_FINAL_COEF_CHECK = "DISABLED";
	parameter SLOT_CLOCK_CONFIGURATION = "REFCLK_BY_SLOT";
	parameter SLOT_IMPLEMENTED = "UNCONNECTED";
	parameter SLOT_POWER_LIMIT_SCALE = "0b00";
	parameter SLOT_POWER_LIMIT_VALUE = "0b00001010";
	parameter SPEED_LPBK_CTRL = "2P5G";
	parameter START_PRESET = "PRESET_VALUE";
	parameter START_REMOTE_ADV = "OTHERWISE";
	parameter STATE_DATA_N = "USE_RX_DATA_OBSERVATION";
	parameter STEP_SELECT = "0b00000";
	parameter STP_OVERRIDE_EN = "DISABLED";
	parameter STP_OVERRIDE_LEN = "0b00000000000";
	parameter STP_OVERRIDE_NEW_LEN = "0b00000000000";
	parameter SUBSTATE_MAX = "0b00000";
	parameter SUBSYSTEM_ID_ID2A = "0b1110000000000100";
	parameter SUBSYSTEM_ID_ID2B = "0b1110000000000100";
	parameter SUBSYSTEM_ID_ID2C = "0b1110000000000100";
	parameter SUBSYSTEM_ID_ID2D = "0b1110000000000100";
	parameter SUBSYSTEM_VENDOR_ID_ID2A = "0b0001100110101010";
	parameter SUBSYSTEM_VENDOR_ID_ID2B = "0b0001100110101010";
	parameter SUBSYSTEM_VENDOR_ID_ID2C = "0b0001100110101010";
	parameter SUBSYSTEM_VENDOR_ID_ID2D = "0b0001100110101010";
	parameter SUPP_SIZE_CFG0_A = "0b00000000000000001111";
	parameter SUPP_SIZE_CFG0_B = "0b00000000000000001111";
	parameter SUPP_SIZE_CFG0_C = "0b00000000000000001111";
	parameter SUPP_SIZE_CFG0_D = "0b00000000000000001111";
	parameter SUPP_SIZE_CFG1_A = "0b00000000000000000000";
	parameter SUPP_SIZE_CFG1_B = "0b00000000000000000000";
	parameter SUPP_SIZE_CFG1_C = "0b00000000000000000000";
	parameter SUPP_SIZE_CFG1_D = "0b00000000000000000000";
	parameter SUPP_SIZE_CFG2_A = "0b00000000000000000000";
	parameter SUPP_SIZE_CFG2_B = "0b00000000000000000000";
	parameter SUPP_SIZE_CFG2_C = "0b00000000000000000000";
	parameter SUPP_SIZE_CFG2_D = "0b00000000000000000000";
	parameter SUPP_SIZE_CFG3_A = "0b00000000000000000000";
	parameter SUPP_SIZE_CFG3_B = "0b00000000000000000000";
	parameter SUPP_SIZE_CFG3_C = "0b00000000000000000000";
	parameter SUPP_SIZE_CFG3_D = "0b00000000000000000000";
	parameter SUPP_SIZE_CFG4_A = "0b00000000000000000000";
	parameter SUPP_SIZE_CFG4_B = "0b00000000000000000000";
	parameter SUPP_SIZE_CFG4_C = "0b00000000000000000000";
	parameter SUPP_SIZE_CFG4_D = "0b00000000000000000000";
	parameter SUPP_SIZE_CFG5_A = "0b00000000000000000000";
	parameter SUPP_SIZE_CFG5_B = "0b00000000000000000000";
	parameter SUPP_SIZE_CFG5_C = "0b00000000000000000000";
	parameter SUPP_SIZE_CFG5_D = "0b00000000000000000000";
	parameter SYS_ALLOC = "PWR_BUDGET_CAP_VALUES";
	parameter T0_RX_BYPASS_MSG_DEC = "NORMAL_OPERATION";
	parameter TABLE_SIZE_MSIXCAP_A = "0b00000000111";
	parameter TABLE_SIZE_MSIXCAP_B = "0b00000000111";
	parameter TABLE_SIZE_MSIXCAP_C = "0b00000000111";
	parameter TABLE_SIZE_MSIXCAP_D = "0b00000000111";
	parameter TARGET_LINK_SPEED = "8G";
	parameter TARGET_ONLY = "DISABLED";
	parameter TD1_MEANS_ADD_HAS_N = "ECRC_CONTAINED";
	parameter TIMEOUT_THRESHOLD_PME = "0b000000000000";
	parameter TIMEOUT_THRESHOLD_PME_TO_ACK_DS = "0b00000000";
	parameter TIMER = "0b00000000";
	parameter TLP_LCRC_ERR_ENABLE = "DISABLED";
	parameter TLP_LCRC_ERR_RATE = "0b000";
	parameter TLP_SEQ_ERR_ENABLE = "DISABLED";
	parameter TLUNIT = "1_MS";
	parameter TO_EXTEND = "0b01111111";
	parameter TRNG_A0COEF = "0b101";
	parameter TRNG_A1COEF = "0b101";
	parameter TRNG_A2COEF = "0b101";
	parameter TRNG_FAST = "DISABLED";
	parameter TRNG_ITERCNT = "0b100";
	parameter TRNG_RXEQ_TIMER = "0b00100000";
	parameter TS1_ACK_BLOCK_USE_PRESET = "FORCED_TO_ZERO";
	parameter TS1_ACK_DELAY = "0b00011111";
	parameter TS1_ACK_MASK_USE_PRESET = "IGNORES_USE_PRESET";
	parameter TX_AMP_RATIO_MARGIN0_FULL = "0b10000000";
	parameter TX_AMP_RATIO_MARGIN0_HALF = "0b01010000";
	parameter TX_AMP_RATIO_MARGIN1_FULL = "0b01111000";
	parameter TX_AMP_RATIO_MARGIN1_HALF = "0b01011000";
	parameter TX_AMP_RATIO_MARGIN2_FULL = "0b01101000";
	parameter TX_AMP_RATIO_MARGIN2_HALF = "0b01001000";
	parameter TX_AMP_RATIO_MARGIN3_FULL = "0b01100000";
	parameter TX_AMP_RATIO_MARGIN3_HALF = "0b01000000";
	parameter TX_AMP_RATIO_MARGIN4_FULL = "0b01011000";
	parameter TX_AMP_RATIO_MARGIN4_HALF = "0b00111000";
	parameter TX_AMP_RATIO_MARGIN5_FULL = "0b01010000";
	parameter TX_AMP_RATIO_MARGIN5_HALF = "0b00110000";
	parameter TX_AMP_RATIO_MARGIN6_FULL = "0b01001000";
	parameter TX_AMP_RATIO_MARGIN6_HALF = "0b00101000";
	parameter TX_AMP_RATIO_MARGIN7_FULL = "0b01000000";
	parameter TX_AMP_RATIO_MARGIN7_HALF = "0b00100000";
	parameter TX_BYPASS_DECODE_EN = "ENABLED";
	parameter TX_BYPASS_MSG_DEC = "NORMAL_OPERATION";
	parameter TX_COMP_RECEIVE = "DOES_NOT_ASSERT";
	parameter TX_CONVERT_UR_TO_CA = "NORMAL_OPERATION";
	parameter TX_D_ALLOC_C = "0b0000000001100000";
	parameter TX_D_ALLOC_N = "0b0000000000000110";
	parameter TX_D_ALLOC_P = "0b0000000001101100";
	parameter TX_DIV_MODE0 = "0b10";
	parameter TX_DIV_MODE1 = "0b10";
	parameter TX_DIV_MODE2 = "0b10";
	parameter TX_EQ_EVAL_CNT_SEL = "WAIT_8_CLKS";
	parameter TX_ERR_COR = "DISABLED";
	parameter TX_ERR_UCOR = "DISABLED";
	parameter TX_FORCE_RO = "DISABLED";
	parameter TX_GAP_INJECT_EN = "DO_NOT_INJECT_GAP";
	parameter TX_H_ALLOC_C = "0b000000100000";
	parameter TX_H_ALLOC_N = "0b000000001000";
	parameter TX_H_ALLOC_P = "0b000000010000";
	parameter TX_HIZ = "IGNORED";
	parameter TX_IMPED_RATIO = "0b10000000";
	parameter TX_PAR1_INJECT_EN = "DO_NOT_INJECT_ERR";
	parameter TX_PAR2_HANDLE_DISABLE = "ENABLE_HANDLING";
	parameter TX_PAR2_INJECT_EN = "DO_NOT_INJECT_ERR";
	parameter TX_PAR2_REPORT_DISABLE = "ENABLE_REPORTING";
	parameter TX_POLINV = "NORMAL";
	parameter TX_PRE_RATIO = "0b00000000";
	parameter TX_PRE_RATIO_DEEMP0_FULL = "0b00000000";
	parameter TX_PRE_RATIO_DEEMP0_HALF = "0b00000000";
	parameter TX_PRE_RATIO_DEEMP1_FULL = "0b00000000";
	parameter TX_PRE_RATIO_DEEMP1_HALF = "0b00000000";
	parameter TX_PRIORITY = "DISABLED";
	parameter TX_PRIORITY_N_STARVE_THRESH = "0b00010000";
	parameter TX_PRIORITY_P_STARVE_THRESH = "0b00010000";
	parameter TX_PST_RATIO = "0b00010101";
	parameter TX_PST_RATIO_DEEMP0_FULL = "0b00100000";
	parameter TX_PST_RATIO_DEEMP0_HALF = "0b00100000";
	parameter TX_PST_RATIO_DEEMP1_FULL = "0b00010101";
	parameter TX_PST_RATIO_DEEMP1_HALF = "0b00010101";
	parameter TX_QUIESCE = "DISABLED";
	parameter TX_REPLAY_ECC1_HANDLE_DISABLE = "ENABLE_CORRECTION";
	parameter TX_REPLAY_ECC1_INJECT_EN = "DO_NOT_INJECT_ERR";
	parameter TX_REPLAY_ECC1_REPORT_DISABLE = "ENABLE_REPORTING";
	parameter TX_REPLAY_ECC2_HANDLE_DISABLE = "ENABLE_HANDLING";
	parameter TX_REPLAY_ECC2_INJECT_EN = "DO_NOT_INJECT_ERR";
	parameter TX_REPLAY_ECC2_REPORT_DISABLE = "ENABLE_REPORTING";
	parameter TX_REQ_EQ = "DISABLED";
	parameter TX_SELECT_RX_FEEDBACK = "REFCLK";
	parameter TX_TLP_VALID = "DISABLED";
	parameter TXF_A = "0b0100";
	parameter TXF_B = "0b0100";
	parameter TXF_C = "0b0100";
	parameter TXHF_CLKDN = "ENABLED";
	parameter TXM_A = "0b10";
	parameter TXM_B = "0b01";
	parameter TXM_C = "0b00";
	parameter TXN_A = "0b00100";
	parameter TXN_B = "0b01001";
	parameter TXN_C = "0b01111";
	parameter TXPLL_INIT = "DISABLED";
	parameter TXPLLRST = "DISABLED";
	parameter TYPE1_TYPE0_N = "ENDPOINT";
	parameter U_CLK_PERIOD = "0b0001111101000000";
	parameter US_PORT_PS_ENTRY_TIME = "0b0000000000000000";
	parameter US_PORT_RX_PRESET_HINT = "0b010";
	parameter US_PORT_TX_PRESET = "0b0100";
	parameter USE_COEF_PRE_MTHD_CTRL = "PRESET_VALUE";
	parameter USE_COEF_UPDN_CTRL = "PRESET_VALUE";
	parameter USER_AUTO_N = "AUTOMATIC_ON_RECEPTION";
	parameter VEC_MASK_CAPABLE_MSICAP_A = "ENABLED";
	parameter VEC_MASK_CAPABLE_MSICAP_B = "ENABLED";
	parameter VEC_MASK_CAPABLE_MSICAP_C = "ENABLED";
	parameter VEC_MASK_CAPABLE_MSICAP_D = "ENABLED";
	parameter VENDOR_ID_ID1A = "0b0001100110101010";
	parameter VENDOR_ID_ID1B = "0b0001100110101010";
	parameter VENDOR_ID_ID1C = "0b0001100110101010";
	parameter VENDOR_ID_ID1D = "0b0001100110101010";
	parameter VENDOR0_UR = "REPORT";
	parameter VERSION_AER_CAP = "VER_0X2";
	parameter VERSION_PM_CAP = "0b011";
	parameter XLCY0 = "0b00000000";
	parameter XLCY1 = "0b00000000";
	parameter RX_ESP_RESP_WAIT = "0b01000000";
	parameter SEL_PCLK_DIV2 = "PCLK_DIV2";
	parameter COMPLIANCE = "ENABLED";
	parameter LOOPBACK = "ENABLED";
	parameter HOT_RESET = "ENABLED";
	parameter DIS_PREVENT = "ENABLED";
	parameter MPS_VIOLATION_RX = "DISABLED";
	parameter MPS_VIOLATION_TX = "DISABLED";
	parameter EN_RX_ALLOC_SEL = "HW";
	parameter EN_TX_ALLOC_SEL = "HW";
	parameter AUX_CLK_PERIOD = "0b1111010000100100";
	parameter EN_PIPE_IF_CTRL = "DISABLED";
	parameter PIPE_PWRDN = "P1";
	parameter TX_CM_DIS = "DEASSERTED";
	parameter RX_EI_DIS = "DEASSERTED";
	parameter PCLKREQ_N = "DEASSERTED";
	parameter STS_PHY_STATUS = "DEASSERTED";
	parameter STS_PIPE_RSTN = "DEASSERTED";
	parameter LEGACY_MODE = "MATCH_TS";
	parameter OVERFLOW = "DISABLED";
	parameter DIR = "RECEIVE";
	parameter SPEED = "8G";
	parameter LANE = "0";
	parameter COEF_ENABLE_8G = "DISABLED";
	parameter PRESET_ENABLE_8G = "DISABLED";
	parameter VALUE_8G_PRE = "0b000000";
	parameter VALUE_8G_POST = "0b000000";
	parameter REQ_EQ_MAX_COUNT = "0b10";
	parameter MESO_LPBK = "DISABLED";
	parameter TX_REPLAY_ECC2_INJECT_M_1_N = "INJECT_1_ERR";
	parameter TX_REPLAY_ECC1_INJECT_M_1_N = "INJECT_1_ERR";
	parameter REDO = "DISABLED";
	parameter RX_PAR_REPORT_DISABLE = "ENABLE_REPORTING";
	parameter RX_PAR_INJECT_EN = "DO_NOT_INJECT_ERR";
	parameter RX_ECC2_REPORT_DISABLE = "ENABLE_REPORTING";
	parameter RX_ECC2_HANDLE_DISABLE = "ENABLE_HANDLING";
	parameter RX_ECC2_INJECT_M_1_N = "INJECT_1_ERR";
	parameter RX_ECC2_INJECT_TYPE = "POSTED_DATA_RAM";
	parameter RX_ECC2_INJECT_EN = "DO_NOT_INJECT_ERR";
	parameter RX_ECC1_REPORT_DISABLE = "ENABLE_REPORTING";
	parameter RX_ECC1_HANDLE_DISABLE = "ENABLE_HANDLING";
	parameter RX_ECC1_INJECT_M_1_N = "INJECT_1_ERR";
	parameter RX_ECC1_INJECT_TYPE = "POSTED_DATA_RAM";
	parameter RX_ECC1_INJECT_EN = "DO_NOT_INJECT_ERR";
	parameter RX_ERR_PAR = "OTHERWISE";
	parameter RX_ERR_ECC2 = "OTHERWISE";
	parameter RX_ERR_ECC1 = "OTHERWISE";
	parameter TX_PAR_REPORT_DISABLE = "ENABLE_REPORTING";
	parameter TX_PAR_INJECT_EN = "DO_NOT_INJECT_ERR";
	parameter TX_ECC2_REPORT_DISABLE = "ENABLE_REPORTING";
	parameter TX_ECC2_HANDLE_DISABLE = "ENABLE_HANDLING";
	parameter TX_ECC2_INJECT_M_1_N = "INJECT_1_ERR";
	parameter TX_ECC2_INJECT_TYPE = "POSTED_DATA_RAM";
	parameter TX_ECC2_INJECT_EN = "DO_NOT_INJECT_ERR";
	parameter TX_ECC1_REPORT_DISABLE = "ENABLE_REPORTING";
	parameter TX_ECC1_HANDLE_DISABLE = "ENABLE_HANDLING";
	parameter TX_ECC1_INJECT_M_1_N = "INJECT_1_ERR";
	parameter TX_ECC1_INJECT_TYPE = "POSTED_DATA_RAM";
	parameter TX_ECC1_INJECT_EN = "DO_NOT_INJECT_ERR";
	parameter TX_ERR_PAR = "OTHERWISE";
	parameter TX_ERR_ECC2 = "OTHERWISE";
	parameter TX_ERR_ECC1 = "OTHERWISE";
	parameter MAX_PAYLOAD_SIZE_SUPPORTED = "256_BYTES";
	parameter ARXCAL_OUT = "DISABLED";
	parameter F_ARXDPDIR = "IGNORED";
	parameter IDLE_INFER_REC_RCVR_CFG = "OTHERWISE";
	parameter IDLE_INFER_LPBK_SLAVE = "OTHERWISE";
	parameter IDLE_INFER_REC_SPEED2_SUCCESS = "OTHERWISE";
	parameter IDLE_INFER_REC_SPEED2_UNSUCCESS = "OTHERWISE";
	parameter IDLE_INFER_L0_TO_REC_RCVR_LOCK = "OTHERWISE";
	parameter SPEED_CHANGE_FAIL = "OTHERWISE";
	parameter DIRECT_TO_DETECT_FAST = "OTHERWISE";
	parameter DIRECT_TO_RCVRY_CH_BOND = "OTHERWISE";
	parameter DIRECT_TO_LPBK_ENTRY = "OTHERWISE";
	parameter DIRECT_SPEED_CHANGE = "OTHERWISE";
	parameter L0_TO_REC_RCVR_LOCK_RX_TS12 = "OTHERWISE";
	parameter L0_TO_REC_RCVR_LOCK_RX_8G_EIE = "OTHERWISE";
	parameter L0_TO_REC_RCVR_LOCK_RX_INFER = "OTHERWISE";
	parameter DIRECT_TO_RCVRY_PHY = "OTHERWISE";
	parameter DIRECT_TO_RCVRY_FRAME = "OTHERWISE";
	parameter DIRECT_TO_RCVRY_REPLAY = "OTHERWISE";
	parameter DIRECT_TO_HOT_RESET = "OTHERWISE";
	parameter DIRECT_TO_DISABLE = "OTHERWISE";
	parameter RX_L0S_DIRECT_TO_RCVRY = "OTHERWISE";
	parameter AUTONOMOUS_WIDTH_CHANGE = "OTHERWISE";
	parameter DIRECTED_RETRAIN_LINK = "OTHERWISE";
	parameter ERR_TX_PIPE_UNDERFLOW = "OTHERWISE";
	parameter TS2_DETECT3 = "OTHERWISE";
	parameter TS2_DETECT2 = "OTHERWISE";
	parameter TS2_DETECT1 = "OTHERWISE";
	parameter TS2_DETECT0 = "OTHERWISE";
	parameter TS1_DETECT3 = "OTHERWISE";
	parameter TS1_DETECT2 = "OTHERWISE";
	parameter TS1_DETECT1 = "OTHERWISE";
	parameter TS1_DETECT0 = "OTHERWISE";
	parameter TS2I_DETECT3 = "OTHERWISE";
	parameter TS2I_DETECT2 = "OTHERWISE";
	parameter TS2I_DETECT1 = "OTHERWISE";
	parameter TS2I_DETECT0 = "OTHERWISE";
	parameter TS1I_DETECT3 = "OTHERWISE";
	parameter TS1I_DETECT2 = "OTHERWISE";
	parameter TS1I_DETECT1 = "OTHERWISE";
	parameter TS1I_DETECT0 = "OTHERWISE";
	parameter FTS_DETECT3 = "OTHERWISE";
	parameter FTS_DETECT2 = "OTHERWISE";
	parameter FTS_DETECT1 = "OTHERWISE";
	parameter FTS_DETECT0 = "OTHERWISE";
	parameter SKP_DETECT3 = "OTHERWISE";
	parameter SKP_DETECT2 = "OTHERWISE";
	parameter SKP_DETECT1 = "OTHERWISE";
	parameter SKP_DETECT0 = "OTHERWISE";
	parameter EIE_DETECT3 = "OTHERWISE";
	parameter EIE_DETECT2 = "OTHERWISE";
	parameter EIE_DETECT1 = "OTHERWISE";
	parameter EIE_DETECT0 = "OTHERWISE";
	parameter EIOS_DETECT3 = "OTHERWISE";
	parameter EIOS_DETECT2 = "OTHERWISE";
	parameter EIOS_DETECT1 = "OTHERWISE";
	parameter EIOS_DETECT0 = "OTHERWISE";
	parameter DATA_DETECT3 = "OTHERWISE";
	parameter DATA_DETECT2 = "OTHERWISE";
	parameter DATA_DETECT1 = "OTHERWISE";
	parameter DATA_DETECT0 = "OTHERWISE";
	parameter SDS_DETECT3 = "OTHERWISE";
	parameter SDS_DETECT2 = "OTHERWISE";
	parameter SDS_DETECT1 = "OTHERWISE";
	parameter SDS_DETECT0 = "OTHERWISE";
	parameter INFO_BAD_TLP_NULL_ERR = "OTHERWISE";
	parameter INFO_BAD_TLP_PHY_ERR = "OTHERWISE";
	parameter INFO_BAD_TLP_MALF_ERR = "OTHERWISE";
	parameter INFO_BAD_TLP_ECRC_ERR = "OTHERWISE";
	parameter INFO_SCHEDULE_DUPL_ACK = "OTHERWISE";
	parameter INFO_BAD_TLP_SEQ_ERR = "OTHERWISE";
	parameter INFO_BAD_TLP_CRC_ERR = "OTHERWISE";
	parameter INFO_NAK_RECEIVED = "OTHERWISE";
	parameter INFO_DESKEW_OVERFLOW_ERROR = "OTHERWISE";
	parameter INFO_TX_DATA_UNDERFLOW = "OTHERWISE";
	parameter INFO_REPLAY_STARTED = "OTHERWISE";
	parameter ERR_AER_TX_PAR2 = "OTHERWISE";
	parameter ERR_AER_TX_REPLAY_ECC2 = "OTHERWISE";
	parameter ERR_AER_TX_REPLAY_ECC1 = "OTHERWISE";
	parameter ERR_AER_SURPRISE_DOWN = "OTHERWISE";
	parameter ERR_AER_DL_PROTOCOL_ERROR = "OTHERWISE";
	parameter ERR_AER_REPLAY_TIMER_TIMEOUT = "OTHERWISE";
	parameter ERR_AER_REPLAY_NUM_ROLLOVER = "OTHERWISE";
	parameter ERR_AER_BAD_DLLP = "OTHERWISE";
	parameter ERR_AER_BAD_TLP = "OTHERWISE";
	parameter ERR_AER_RECEIVER_ERROR = "OTHERWISE";
	parameter P_RX_LIM_H = "DISABLED";
	parameter P_RX_LIM_D = "DISABLED";
	parameter N_RX_LIM_H = "DISABLED";
	parameter N_RX_LIM_D = "DISABLED";
	parameter C_RX_LIM_H = "DISABLED";
	parameter C_RX_LIM_D = "DISABLED";
	parameter P_TX_LIM_H = "DISABLED";
	parameter P_TX_LIM_D = "DISABLED";
	parameter N_TX_LIM_H = "DISABLED";
	parameter N_TX_LIM_D = "DISABLED";
	parameter C_TX_LIM_H = "DISABLED";
	parameter C_TX_LIM_D = "DISABLED";
	parameter MAX_RSA_WAIT = "0b00101000";
	parameter F_ARXDPNULL = "0b00000";

endmodule


module PLL_CORE (CIBDIR, CIBDSEL2, CIBDSEL1, CIBDSEL0, CIBLDREG, CIBROT, CLKOP, CLKOS, CLKOS2, CLKOS3, CLKOS4, CLKOS5, ENEXT, ENCLKOP, ENCLKOS, ENCLKOS2, ENCLKOS3, ENCLKOS4, ENCLKOS5, FBKCK, INTFBK5, INTFBK4, INTFBK3, INTFBK2, INTFBK1, INTFBK0, INTLOCK, LEGACY, LEGRDYN, LMMICLK, LMMIOFFSET6, LMMIOFFSET5, LMMIOFFSET4, LMMIOFFSET3, LMMIOFFSET2, LMMIOFFSET1, LMMIOFFSET0, LMMIRDATA7, LMMIRDATA6, LMMIRDATA5, LMMIRDATA4, LMMIRDATA3, LMMIRDATA2, LMMIRDATA1, LMMIRDATA0, LMMIRDATAVALID, LMMIREADY, LMMIREQUEST, LMMIRESETN, LMMIWDATA7, LMMIWDATA6, LMMIWDATA5, LMMIWDATA4, LMMIWDATA3, LMMIWDATA2, LMMIWDATA1, LMMIWDATA0, LMMIWRRDN, LOCK, PFDDN, PFDUP, PLLRESET, REFCK, STDBY, ZRSEL3, REFMUXCK, PLLPDN, REGQA, REGQB, REGQB1, CLKOUTDL, ROTDEL, DIRDEL, ROTDELP1, GRAYTEST4, GRAYTEST3, GRAYTEST2, GRAYTEST1, GRAYTEST0, BINTEST1, BINTEST0, DIRDELP1, GRAYACT4, GRAYACT3, GRAYACT2, GRAYACT1, GRAYACT0, BINACT1, BINACT0, OPCGLDCK, SCANRST, SCANCLK, REFDETRESET, REFDETLOS); //synthesis syn_black_box syn_lib_cell=1

	input CIBDIR;
	input CIBDSEL2;
	input CIBDSEL1;
	input CIBDSEL0;
	input CIBLDREG;
	input CIBROT;
	output CLKOP;
	output CLKOS;
	output CLKOS2;
	output CLKOS3;
	output CLKOS4;
	output CLKOS5;
	input ENEXT;
	input ENCLKOP;
	input ENCLKOS;
	input ENCLKOS2;
	input ENCLKOS3;
	input ENCLKOS4;
	input ENCLKOS5;
	input FBKCK;
	output INTFBK5;
	output INTFBK4;
	output INTFBK3;
	output INTFBK2;
	output INTFBK1;
	output INTFBK0;
	output INTLOCK;
	input LEGACY;
	output LEGRDYN;
	input LMMICLK;
	input LMMIOFFSET6;
	input LMMIOFFSET5;
	input LMMIOFFSET4;
	input LMMIOFFSET3;
	input LMMIOFFSET2;
	input LMMIOFFSET1;
	input LMMIOFFSET0;
	output LMMIRDATA7;
	output LMMIRDATA6;
	output LMMIRDATA5;
	output LMMIRDATA4;
	output LMMIRDATA3;
	output LMMIRDATA2;
	output LMMIRDATA1;
	output LMMIRDATA0;
	output LMMIRDATAVALID;
	output LMMIREADY;
	input LMMIREQUEST;
	input LMMIRESETN;
	input LMMIWDATA7;
	input LMMIWDATA6;
	input LMMIWDATA5;
	input LMMIWDATA4;
	input LMMIWDATA3;
	input LMMIWDATA2;
	input LMMIWDATA1;
	input LMMIWDATA0;
	input LMMIWRRDN;
	output LOCK;
	output PFDDN;
	output PFDUP;
	input PLLRESET;
	input REFCK;
	input STDBY;
	input ZRSEL3;
	output REFMUXCK;
	input PLLPDN;
	output REGQA;
	output REGQB;
	output REGQB1;
	output CLKOUTDL;
	input ROTDEL;
	input DIRDEL;
	input ROTDELP1;
	input GRAYTEST4;
	input GRAYTEST3;
	input GRAYTEST2;
	input GRAYTEST1;
	input GRAYTEST0;
	input BINTEST1;
	input BINTEST0;
	input DIRDELP1;
	input GRAYACT4;
	input GRAYACT3;
	input GRAYACT2;
	input GRAYACT1;
	input GRAYACT0;
	input BINACT1;
	input BINACT0;
	input OPCGLDCK;
	input SCANRST;
	input SCANCLK;
	input REFDETRESET;
	output REFDETLOS;

	parameter BW_CTL_BIAS = "0b0101";
	parameter CLKOP_TRIM = "0b0000";
	parameter CLKOS_TRIM = "0b0000";
	parameter CLKOS2_TRIM = "0b0000";
	parameter CLKOS3_TRIM = "0b0000";
	parameter CLKOS4_TRIM = "0b0000";
	parameter CLKOS5_TRIM = "0b0000";
	parameter CRIPPLE = "5P";
	parameter CSET = "40P";
	parameter DELAY_CTRL = "200PS";
	parameter DELA = "0";
	parameter DELB = "0";
	parameter DELC = "0";
	parameter DELD = "0";
	parameter DELE = "0";
	parameter DELF = "0";
	parameter DIRECTION = "DISABLED";
	parameter DIVA = "0";
	parameter DIVB = "0";
	parameter DIVC = "0";
	parameter DIVD = "0";
	parameter DIVE = "0";
	parameter DIVF = "0";
	parameter DYN_SEL = "0b000";
	parameter DYN_SOURCE = "STATIC";
	parameter ENCLK_CLKOP = "DISABLED";
	parameter ENCLK_CLKOS = "DISABLED";
	parameter ENCLK_CLKOS2 = "DISABLED";
	parameter ENCLK_CLKOS3 = "DISABLED";
	parameter ENCLK_CLKOS4 = "DISABLED";
	parameter ENCLK_CLKOS5 = "DISABLED";
	parameter ENABLE_SYNC = "DISABLED";
	parameter FAST_LOCK_EN = "ENABLED";
	parameter V2I_1V_EN = "DISABLED";
	parameter FBK_CUR_BLE = "0b00000000";
	parameter FBK_EDGE_SEL = "POSITIVE";
	parameter FBK_IF_TIMING_CTL = "0b00";
	parameter FBK_INTEGER_MODE = "DISABLED";
	parameter FBK_MASK = "0b00001000";
	parameter FBK_MMD_DIG = "8";
	parameter FBK_MMD_PULS_CTL = "0b0000";
	parameter FBK_MODE = "0b00";
	parameter FBK_PI_BYPASS = "NOT_BYPASSED";
	parameter FBK_PI_RC = "0b1100";
	parameter FBK_PR_CC = "0b0000";
	parameter FBK_PR_IC = "0b1000";
	parameter FLOAT_CP = "DISABLED";
	parameter FLOCK_CTRL = "2X";
	parameter FLOCK_EN = "ENABLED";
	parameter FLOCK_SRC_SEL = "REFCLK";
	parameter FORCE_FILTER = "DISABLED";
	parameter I_CTRL = "10UA";
	parameter IPI_CMP = "0b1000";
	parameter IPI_CMPN = "0b0011";
	parameter IPI_COMP_EN = "DISABLED";
	parameter IPP_CTRL = "0b1000";
	parameter IPP_SEL = "0b1111";
	parameter KP_VCO = "0b11001";
	parameter LDT_INT_LOCK_STICKY = "DISABLED";
	parameter LDT_LOCK = "1536CYC";
	parameter LDT_LOCK_SEL = "U_FREQ";
	parameter LEGACY_ATT = "DISABLED";
	parameter LOAD_REG = "DISABLED";
	parameter OPENLOOP_EN = "DISABLED";
	parameter PHIA = "0";
	parameter PHIB = "0";
	parameter PHIC = "0";
	parameter PHID = "0";
	parameter PHIE = "0";
	parameter PHIF = "0";
	parameter PLLPDN_EN = "DISABLED";
	parameter PLLPD_N = "UNUSED";
	parameter PLLRESET_ENA = "DISABLED";
	parameter REF_INTEGER_MODE = "DISABLED";
	parameter REF_MASK = "0b00000000";
	parameter REF_MMD_DIG = "8";
	parameter REF_MMD_IN = "0b00001000";
	parameter REF_MMD_PULS_CTL = "0b0000";
	parameter REF_TIMING_CTL = "0b00";
	parameter REFIN_RESET = "SET";
	parameter RESET_LF = "DISABLED";
	parameter ROTATE = "DISABLED";
	parameter SEL_OUTA = "DISABLED";
	parameter SEL_OUTB = "DISABLED";
	parameter SEL_OUTC = "DISABLED";
	parameter SEL_OUTD = "DISABLED";
	parameter SEL_OUTE = "DISABLED";
	parameter SEL_OUTF = "DISABLED";
	parameter SLEEP = "DISABLED";
	parameter SSC_DITHER = "DISABLED";
	parameter SSC_EN_CENTER_IN = "DOWN_TRIANGLE";
	parameter SSC_EN_SDM = "DISABLED";
	parameter SSC_EN_SSC = "DISABLED";
	parameter SSC_F_CODE = "0b000000000000000";
	parameter SSC_N_CODE = "0b000010100";
	parameter SSC_ORDER = "SDM_ORDER2";
	parameter SSC_PI_BYPASS = "NOT_BYPASSED";
	parameter SSC_REG_WEIGHTING_SEL = "0b000";
	parameter SSC_SQUARE_MODE = "DISABLED";
	parameter SSC_STEP_IN = "0b0000000";
	parameter SSC_TBASE = "0b000000000000";
	parameter STDBY_ATT = "DISABLED";
	parameter TRIMOP_BYPASS_N = "BYPASSED";
	parameter TRIMOS_BYPASS_N = "BYPASSED";
	parameter TRIMOS2_BYPASS_N = "BYPASSED";
	parameter TRIMOS3_BYPASS_N = "BYPASSED";
	parameter TRIMOS4_BYPASS_N = "BYPASSED";
	parameter TRIMOS5_BYPASS_N = "BYPASSED";
	parameter V2I_KVCO_SEL = "85";
	parameter V2I_PP_ICTRL = "0b00110";
	parameter V2I_PP_RES = "10K";
	parameter CLKMUX_FB = "CMUX_CLKOP";
	parameter SEL_FBK = "DIVA";
	parameter DIV_DEL = "0b0000001";
	parameter PHASE_SEL_DEL = "0b000";
	parameter PHASE_SEL_DEL_P1 = "0b000";
	parameter EXTERNAL_DIVIDE_FACTOR = "0";
	parameter INTFBKDEL_SEL = "DISABLED";
	parameter PMU_WAITFORLOCK = "ENABLED";
	parameter REF_OSC_CTRL = "3P2";
	parameter REF_COUNTS = "0000";
	parameter REF_USE = "DISABLED";
	parameter REF_ENABLE = "DISABLED";
	parameter SIM_FLOAT_PRECISION = "0.0001";

endmodule


module PREADD9_CORE (B8, B7, B6, B5, B4, B3, B2, B1, B0, BSIGNED, C9, C8, C7, C6, C5, C4, C3, C2, C1, C0, BRS18, BRS17, BRS16, BRS15, BRS14, BRS13, BRS12, BRS11, BRS10, BRS28, BRS27, BRS26, BRS25, BRS24, BRS23, BRS22, BRS21, BRS20, BLS18, BLS17, BLS16, BLS15, BLS14, BLS13, BLS12, BLS11, BLS10, BLS28, BLS27, BLS26, BLS25, BLS24, BLS23, BLS22, BLS21, BLS20, BRSS1, BRSS2, BLSS1, BLSS2, PRCASIN, CLK, RSTB, CEB, RSTCL, CECL, BRSO8, BRSO7, BRSO6, BRSO5, BRSO4, BRSO3, BRSO2, BRSO1, BRSO0, BLSO8, BLSO7, BLSO6, BLSO5, BLSO4, BLSO3, BLSO2, BLSO1, BLSO0, BRSOSGND, BLSOSGND, PRCASOUT, BR8, BR7, BR6, BR5, BR4, BR3, BR2, BR1, BR0, BRSIGNED); //synthesis syn_black_box syn_lib_cell=1

	input B8;
	input B7;
	input B6;
	input B5;
	input B4;
	input B3;
	input B2;
	input B1;
	input B0;
	input BSIGNED;
	input C9;
	input C8;
	input C7;
	input C6;
	input C5;
	input C4;
	input C3;
	input C2;
	input C1;
	input C0;
	input BRS18;
	input BRS17;
	input BRS16;
	input BRS15;
	input BRS14;
	input BRS13;
	input BRS12;
	input BRS11;
	input BRS10;
	input BRS28;
	input BRS27;
	input BRS26;
	input BRS25;
	input BRS24;
	input BRS23;
	input BRS22;
	input BRS21;
	input BRS20;
	input BLS18;
	input BLS17;
	input BLS16;
	input BLS15;
	input BLS14;
	input BLS13;
	input BLS12;
	input BLS11;
	input BLS10;
	input BLS28;
	input BLS27;
	input BLS26;
	input BLS25;
	input BLS24;
	input BLS23;
	input BLS22;
	input BLS21;
	input BLS20;
	input BRSS1;
	input BRSS2;
	input BLSS1;
	input BLSS2;
	input PRCASIN;
	input CLK;
	input RSTB;
	input CEB;
	input RSTCL;
	input CECL;
	output BRSO8;
	output BRSO7;
	output BRSO6;
	output BRSO5;
	output BRSO4;
	output BRSO3;
	output BRSO2;
	output BRSO1;
	output BRSO0;
	output BLSO8;
	output BLSO7;
	output BLSO6;
	output BLSO5;
	output BLSO4;
	output BLSO3;
	output BLSO2;
	output BLSO1;
	output BLSO0;
	output BRSOSGND;
	output BLSOSGND;
	output PRCASOUT;
	output BR8;
	output BR7;
	output BR6;
	output BR5;
	output BR4;
	output BR3;
	output BR2;
	output BR1;
	output BR0;
	output BRSIGNED;

	parameter SIGNEDSTATIC_EN = "DISABLED";
	parameter SUBSTRACT_EN = "SUBTRACTION";
	parameter CSIGNED = "DISABLED";
	parameter BSIGNED_OPERAND_EN = "DISABLED";
	parameter BYPASS_PREADD9 = "USED";
	parameter REGBYPSBR0 = "REGISTER";
	parameter REGBYPSBR1 = "BYPASS";
	parameter REGBYPSBL = "REGISTER";
	parameter SHIFTBR = "REGISTER";
	parameter SHIFTBL = "REGISTER";
	parameter GSR = "ENABLED";
	parameter PREADDCAS_EN = "DISABLED";
	parameter SR_18BITSHIFT_EN = "DISABLED";
	parameter OPC = "INPUT_B_AS_PREADDER_OPERAND";
	parameter RESET = "SYNC";

endmodule

module REFMUX_CORE (REFCK, ZRSEL3, REFSEL, REFCLK17, REFCLK16, REFCLK15, REFCLK14, REFCLK13, REFCLK12, REFCLK11, REFCLK10, REFCLK27, REFCLK26, REFCLK25, REFCLK24, REFCLK23, REFCLK22, REFCLK21, REFCLK20); //synthesis syn_black_box syn_lib_cell=1

	output REFCK;
	output ZRSEL3;
	input REFSEL;
	input REFCLK17;
	input REFCLK16;
	input REFCLK15;
	input REFCLK14;
	input REFCLK13;
	input REFCLK12;
	input REFCLK11;
	input REFCLK10;
	input REFCLK27;
	input REFCLK26;
	input REFCLK25;
	input REFCLK24;
	input REFCLK23;
	input REFCLK22;
	input REFCLK21;
	input REFCLK20;

	parameter REFSEL_ATT = "MC1";
	parameter SEL1 = "SELECT_REFCLK1";
	parameter SEL_REF2 = "REFCLK2_0";
	parameter SEL_REF1 = "REFCLK1_0";

endmodule

module REG18_CORE (PM17, PM16, PM15, PM14, PM13, PM12, PM11, PM10, PM9, PM8, PM7, PM6, PM5, PM4, PM3, PM2, PM1, PM0, PP17, PP16, PP15, PP14, PP13, PP12, PP11, PP10, PP9, PP8, PP7, PP6, PP5, PP4, PP3, PP2, PP1, PP0, CEP, RSTP, CLK); //synthesis syn_black_box syn_lib_cell=1

	input PM17;
	input PM16;
	input PM15;
	input PM14;
	input PM13;
	input PM12;
	input PM11;
	input PM10;
	input PM9;
	input PM8;
	input PM7;
	input PM6;
	input PM5;
	input PM4;
	input PM3;
	input PM2;
	input PM1;
	input PM0;
	output PP17;
	output PP16;
	output PP15;
	output PP14;
	output PP13;
	output PP12;
	output PP11;
	output PP10;
	output PP9;
	output PP8;
	output PP7;
	output PP6;
	output PP5;
	output PP4;
	output PP3;
	output PP2;
	output PP1;
	output PP0;
	input CEP;
	input RSTP;
	input CLK;

	parameter REGBYPS = "REGISTER";
	parameter GSR = "ENABLED";
	parameter RESET = "SYNC";

endmodule

module SEIO18_CORE (I, DOLP, B, O, INLP, T, INADC); //synthesis syn_black_box black_box_pad_pin="B" syn_lib_cell=1

	input I;
	input DOLP;
	inout B;
	output O;
	output INLP;
	input T;
	output INADC;

	parameter MIPI_ID = "0";
	parameter PULLMODE = "DOWN";
	parameter MIPI = "DISABLED";
	parameter ENADC_IN = "DISABLED";

endmodule

module SEIO33_CORE (B, O, I, T, I3CRESEN, I3CWKPU); //synthesis syn_black_box black_box_pad_pin="B" syn_lib_cell=1

	inout B;
	output O;
	input I;
	input T;
	input I3CRESEN;
	input I3CWKPU;

	parameter PULLMODE = "DOWN";

endmodule

module SGMIICDR_CORE (DCALIRST, DFACQRST, RRST, SPCLK, SRCLK, SRXD9, SRXD8, SRXD7, SRXD6, SRXD5, SRXD4, SRXD3, SRXD2, SRXD1, SRXD0, LMMICLK, LMMIREQUEST, LMMIWRRDN, LMMIOFFSET3, LMMIOFFSET2, LMMIOFFSET1, LMMIOFFSET0, LMMIWDATA7, LMMIWDATA6, LMMIWDATA5, LMMIWDATA4, LMMIWDATA3, LMMIWDATA2, LMMIWDATA1, LMMIWDATA0, LMMIRDATA7, LMMIRDATA6, LMMIRDATA5, LMMIRDATA4, LMMIRDATA3, LMMIRDATA2, LMMIRDATA1, LMMIRDATA0, LMMIRDATAVALID, LMMIREADY, LMMIRESETN, RSTBFBW, RSTBRXF, SGMIIIN, SREFCLK, CDRLOL, OPCGLOADCLK, SCANCLK, SCANRST); //synthesis syn_black_box syn_lib_cell=1

	input DCALIRST;
	input DFACQRST;
	input RRST;
	input SPCLK;
	output SRCLK;
	output SRXD9;
	output SRXD8;
	output SRXD7;
	output SRXD6;
	output SRXD5;
	output SRXD4;
	output SRXD3;
	output SRXD2;
	output SRXD1;
	output SRXD0;
	input LMMICLK;
	input LMMIREQUEST;
	input LMMIWRRDN;
	input LMMIOFFSET3;
	input LMMIOFFSET2;
	input LMMIOFFSET1;
	input LMMIOFFSET0;
	input LMMIWDATA7;
	input LMMIWDATA6;
	input LMMIWDATA5;
	input LMMIWDATA4;
	input LMMIWDATA3;
	input LMMIWDATA2;
	input LMMIWDATA1;
	input LMMIWDATA0;
	output LMMIRDATA7;
	output LMMIRDATA6;
	output LMMIRDATA5;
	output LMMIRDATA4;
	output LMMIRDATA3;
	output LMMIRDATA2;
	output LMMIRDATA1;
	output LMMIRDATA0;
	output LMMIRDATAVALID;
	output LMMIREADY;
	input LMMIRESETN;
	input RSTBFBW;
	input RSTBRXF;
	input SGMIIIN;
	input SREFCLK;
	output CDRLOL;
	input OPCGLOADCLK;
	input SCANCLK;
	input SCANRST;

	parameter GSR = "ENABLED";
	parameter DCOITUNE4LSB = "0_PERCENT";
	parameter DCOCTLGI = "60_PERCENT";
	parameter DCOSTEP = "17_PERCENT";
	parameter DCOCALDIV = "100_PERCENT";
	parameter DCOIOSTUNE = "49_PERCENT";
	parameter DCOFLTDAC = "181MHZ";
	parameter DCOSTARTVAL = "100_PERCENT";
	parameter DCONUOFLSB = "60_PERCENT";
	parameter RPWDNB = "POWER_UP";
	parameter CDR_CNT4SEL = "BY_4";
	parameter DCOITUNE = "100_PERCENT";
	parameter BAND_THRESHOLD = "0b000000";
	parameter AUTO_FACQ_EN = "ENABLED";
	parameter AUTO_CALIB_EN = "ENABLED";
	parameter CDR_LOL_SET = "2000_PPM";
	parameter FC2DCO_FLOOP = "DISABLED";
	parameter FC2DCO_DLOOP = "DISABLED";
	parameter CALIB_TIME_SEL = "24_CYC";
	parameter CALIB_CK_MODE = "BY_2";
	parameter BAND_CALIB_MODE = "256_FDBK_CLK_CYC";
	parameter REG_BAND_SEL = "0b10101";
	parameter REG_BAND_OFFSET = "0b0000";
	parameter REG_IDAC_SEL = "0b10000000";
	parameter LB_CTL = "DISABLED";
	parameter REG_IDAC_EN = "DISABLED";
	parameter ATDCFG = "0_PS";
	parameter ATDDLY = "0_PS";
	parameter BDAVOID_ENB = "ENABLED";
	parameter BYPASSATD = "NOT_BYPASS";
	parameter DCOIUPDNX2 = "2X";
	parameter IDAC_EN = "DISABLED";
	parameter FB_CLK_DIV = "0b010";
	parameter EN_RECALIB = "ENABLED";

endmodule

module SLICEREG(DL, DF, CLK, LSR, CE, Q); // synthesis syn_black_box syn_lib_cell=1
	input DL;
	input DF;
	input CLK;
	input LSR;
	input CE;
	output Q;
	parameter SEL = "DL";
	parameter REGSET = "RESET";
	parameter LSRMODE = "LSR";
    parameter GSR = "ENABLED";
    parameter ASYNC = "YES";
endmodule


module LUT4(A, B, C, D, Z); // synthesis syn_black_box syn_lib_cell=1
	input A;
	input B;
	input C;
	input D;
	output Z;
	parameter INIT = "0x0000";
endmodule


module SLICEMUX(D1, D0, SEL, Z); // synthesis syn_black_box syn_lib_cell=1
	input D1;
	input D0;
	input SEL;
	output Z;
endmodule


module CCU2(A1, B1, C1, D1, A0, B0, C0, D0, CIN, COUT, S1, S0); // synthesis syn_black_box syn_unconnected_inputs = "CIN" syn_lib_cell=1
	input A1;
	input B1;
	input C1;
	input D1;
	input A0;
	input B0;
	input C0;
	input D0;
	input CIN;
	output COUT;
	output S1;
	output S0;
	parameter INJECT = "YES";
	parameter INIT0 = "0x0000";
	parameter INIT1 = "0x1111";
endmodule


module DPRAM(RAD0, RAD1, RAD2, RAD3, DI0, DI1, WAD0, WAD1, WAD2, WAD3, WCK, WRE, DO1, DO0); // synthesis syn_black_box syn_lib_cell=1
	input RAD0;
	input RAD1;
	input RAD2;
	input RAD3;
	input DI0;
	input DI1;
	input WAD0;
	input WAD1;
	input WAD2;
	input WAD3;
	input WCK;
	input WRE;
	output DO1;
	output DO0;
	parameter INIT0 = "0x0000";
	parameter INIT1 = "0x0000";
endmodule


module IB(I, O); // synthesis syn_black_box black_box_pad_pin="I" syn_lib_cell=1
    input I;
    output O;
endmodule

module OB(I, O); // synthesis syn_black_box black_box_pad_pin="O" syn_lib_cell=1
    input I;
    output O;
endmodule

module OBZ(I, T, O); // synthesis syn_black_box black_box_pad_pin="O" syn_lib_cell=1
    input I;
    input T;
    output O;
endmodule

module FD1P3BX(D, CK, SP, PD, Q); // synthesis syn_black_box syn_lib_cell=1
    input D;
    input CK;
    input SP;
    input PD;
    output Q;
    parameter GSR = "ENABLED";
endmodule

module FD1P3DX(D, CK, SP, CD, Q); // synthesis syn_black_box syn_lib_cell=1
    input D;
    input CK;
    input SP;
    input CD;
    output Q;
    parameter GSR = "ENABLED";
endmodule

module FD1P3IX(D, CK, SP, CD, Q); // synthesis syn_black_box syn_lib_cell=1
    input D;
    input CK;
    input SP;
    input CD;
    output Q;
    parameter GSR = "ENABLED";
endmodule

module FD1P3JX(D, CK, SP, PD, Q); // synthesis syn_black_box syn_lib_cell=1
    input D;
    input CK;
    input SP;
    input PD;
    output Q;
    parameter GSR = "ENABLED";
endmodule

module WIDEFN9(A0, B0, C0, D0, A1, B1, C1, D1, SEL, Z); // synthesis syn_black_box syn_lib_cell=1
    input A0;
    input B0;
    input C0;
    input D0;
    input A1;
    input B1;
    input C1;
    input D1;
    input SEL;
    output Z;
    parameter INIT0 = "0x0000";
    parameter INIT1 = "0x0000";
endmodule

module DPR16X4(RAD, DI, WAD, WRE, WCK, DO); // synthesis syn_black_box syn_lib_cell=1
    input [3:0] RAD;
    input [3:0] DI;
    input [3:0] WAD;
    input WRE;
    input WCK;
    output [3:0] DO;
    parameter INITVAL = "0x0000000000000000";
endmodule

module SPR16X4(DI, CK, WRE, AD, DO); // synthesis syn_black_box syn_lib_cell=1
    input [3:0] DI;
    input CK;
    input WRE;
    input [3:0] AD;
    output [3:0] DO;
    parameter INITVAL = "0x0000000000000000";
endmodule

module GSR(GSR_N, CLK); //synthesis syn_black_box syn_lib_cell=1 syn_noprune=1
    input GSR_N;
    input CLK;
    parameter SYNCMODE = "ASYNC";
endmodule

module DCC (CE, CLKI, CLKO); //synthesis syn_black_box syn_lib_cell=1

	input CE;
	input CLKI;
	output CLKO;

	parameter DCCEN = "0";

endmodule

module DCS (CLK0, CLK1, DCSOUT, SEL, SELFORCE); //synthesis syn_black_box syn_lib_cell=1

	input CLK0;
	input CLK1;
	output DCSOUT;
	input SEL;
	input SELFORCE;

	parameter DCSMODE = "GND";

endmodule

module GSR_CORE (GSROUT, CLK, GSR_N); //synthesis syn_black_box syn_lib_cell=1 syn_noprune=1

	output GSROUT;
	input CLK;
	input GSR_N;

	parameter GSR = "ENABLED";
	parameter GSR_SYNC = "ASYNC";

endmodule

module PCLKDIV (CLKIN, CLKOUT, LSRPDIV, PCLKDIVTESTINP2, PCLKDIVTESTINP1, PCLKDIVTESTINP0); //synthesis syn_black_box syn_lib_cell=1

	input CLKIN;
	output CLKOUT;
	input LSRPDIV;
	input PCLKDIVTESTINP2;
	input PCLKDIVTESTINP1;
	input PCLKDIVTESTINP0;

	parameter DIV_PCLKDIV = "X1";
	parameter GSR = "ENABLED";
	parameter TESTEN_PCLKDIV = "0";
	parameter TESTMODE_PCLKDIV = "0";

endmodule

module VHI (Z); //synthesis syn_black_box syn_lib_cell=1

	output Z;


endmodule

module BB (T, I, O, B); //synthesis syn_black_box black_box_pad_pin="B" syn_lib_cell=1
	input T;
	input I;
	output O;
	inout B;

endmodule

module VLO (Z);  //synthesis syn_black_box syn_lib_cell=1
   output Z ;
endmodule

module INV (A, Z);  //synthesis syn_black_box syn_lib_cell=1
   input A;
   output Z;
endmodule

module BUF (A, Z);  //synthesis syn_black_box syn_lib_cell=1
   input A;
   output Z;
endmodule

module PUR (PUR); // synthesis syn_black_box syn_lib_cell=1 syn_noprune=1
  input PUR;
  parameter RST_PULSE = "1";
endmodule

module RAMW(WD3, WD2, WD1, WD0, WAD3, WAD2, WAD1, WAD0, WCK, WRE, WDO3, WDO2, WDO1, WDO0, WADO3, WADO2, WADO1, WADO0, WCKO, WREO); // synthesis syn_black_box syn_lib_cell=1
    input WD3;
    input WD2;
    input WD1;
    input WD0;
    input WAD3;
    input WAD2;
    input WAD1;
    input WAD0;
    input WCK;
    input WRE;
    output WDO3;
    output WDO2;
    output WDO1;
    output WDO0;
    output WADO3;
    output WADO2;
    output WADO1;
    output WADO0;
    output WCKO;
    output WREO;
endmodule

module IOREG(D, CE, LSR, CLK, Q); // synthesis syn_black_box syn_lib_cell=1
    input D;
    input CE;
    input LSR;
    input CLK;
    output Q;
    parameter REGSET = "RESET";
    parameter ASYNC = "YES";
    parameter GSR = "ENABLED";
endmodule

module PCLKDIVSP(CLKIN, CLKOUT, LSRPDIV); // synthesis syn_black_box syn_lib_cell=1
    input CLKIN;
    output CLKOUT;
    input LSRPDIV;
    parameter DIV_PCLKDIV = "X1";
    parameter GSR = "ENABLED";
endmodule

module JTAGH19 (TDI, TCK, TMS, TDO, JTCK, JTDI, JSHIFT, JUPDATE, JRSTN, JCE2, CDN, IP_ENABLE, ER2_TDO); //synthesis syn_black_box black_box_pad_pin="TDI,TCK,TMS,TDO" syn_lib_cell=1
  input TDI;
  input TCK;
  output TDO;
  input TMS;
  output JTCK;
  output JTDI;
  output JSHIFT;
  output JUPDATE;
  output JRSTN;
  output JCE2;
  output CDN;
  output [18:0] IP_ENABLE;
  input [18:0] ER2_TDO;

  parameter LSCC_FAMILY = "JEDI";
  parameter JTAGHUB_ID = "0x43";
  parameter IP_ENABLE_VAL = "0x00000";
  parameter HUB_00 = "0b0";
  parameter HUB_01 = "0b0";
  parameter HUB_02 = "0b0";
  parameter HUB_03 = "0b0";
  parameter HUB_04 = "0b0";
  parameter HUB_05 = "0b0";
  parameter HUB_06 = "0b0";
  parameter HUB_07 = "0b0";
  parameter HUB_08 = "0b0";
  parameter HUB_09 = "0b0";
  parameter HUB_10 = "0b0";
  parameter HUB_11 = "0b0";
  parameter HUB_12 = "0b0";
  parameter HUB_13 = "0b0";
  parameter HUB_14 = "0b0";
  parameter HUB_15 = "0b0";
  parameter HUB_16 = "0b0";
  parameter HUB_17 = "0b0";
  parameter HUB_18 = "0b0";
endmodule

module JTAGH19SOFT (TDI, TCK, TMS, TDO, JTCK, JTDI, JSHIFT, JUPDATE, JRSTN, JCE2, CDN, IP_ENABLE, ER2_TDO); //synthesis syn_black_box black_box_pad_pin="TDI,TCK,TMS,TDO" syn_lib_cell=1
  input TDI;
  input TCK;
  output TDO;
  input TMS;
  output JTCK;
  output JTDI;
  output JSHIFT;
  output JUPDATE;
  output JRSTN;
  output JCE2;
  output CDN;
  output [18:0] IP_ENABLE;
  input [18:0] ER2_TDO;

  parameter LSCC_FAMILY = "JEDI";
  parameter JTAGHUB_ID = "0x43";
  parameter IP_ENABLE_VAL = "0x00000";
  parameter HUB_00 = "0b0";
  parameter HUB_01 = "0b0";
  parameter HUB_02 = "0b0";
  parameter HUB_03 = "0b0";
  parameter HUB_04 = "0b0";
  parameter HUB_05 = "0b0";
  parameter HUB_06 = "0b0";
  parameter HUB_07 = "0b0";
  parameter HUB_08 = "0b0";
  parameter HUB_09 = "0b0";
  parameter HUB_10 = "0b0";
  parameter HUB_11 = "0b0";
  parameter HUB_12 = "0b0";
  parameter HUB_13 = "0b0";
  parameter HUB_14 = "0b0";
  parameter HUB_15 = "0b0";
  parameter HUB_16 = "0b0";
  parameter HUB_17 = "0b0";
  parameter HUB_18 = "0b0";
endmodule
