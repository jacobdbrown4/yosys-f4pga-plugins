(* top =  1  *)
module lattice_crosslink_nx_evn(gsrn, serial_rx, serial_tx, user_led0, user_led1, user_led2, user_led3, user_led4, user_led5, user_led6, user_led7, user_led8, user_led9, user_led10, user_led11, user_led12, user_led13);
  (* src = "lattice_riscv.v:50640.6-50640.11" *)
  wire CLKOS;
  (* src = "lattice_riscv.v:50641.6-50641.12" *)
  wire CLKOS2;
  (* src = "lattice_riscv.v:50642.6-50642.12" *)
  wire CLKOS3;
  (* src = "lattice_riscv.v:50643.6-50643.12" *)
  wire CLKOS4;
  (* src = "lattice_riscv.v:50652.6-50652.14" *)
  wire CLKOUTDL;
  (* src = "lattice_riscv.v:50693.6-50693.11" *)
  wire CO0_0_TMR_0;
  (* src = "lattice_riscv.v:50693.6-50693.11" *)
  wire CO0_0_TMR_1;
  (* src = "lattice_riscv.v:50693.6-50693.11" *)
  wire CO0_0_TMR_2;
  (* src = "lattice_riscv.v:50692.6-50692.9" *)
  wire CO0_TMR_0;
  (* src = "lattice_riscv.v:50692.6-50692.9" *)
  wire CO0_TMR_1;
  (* src = "lattice_riscv.v:50692.6-50692.9" *)
  wire CO0_TMR_2;
  (* src = "lattice_riscv.v:50724.6-50724.18" *)
  wire FD1P3BX_1_QN;
  (* src = "lattice_riscv.v:50723.6-50723.18" *)
  wire FD1P3BX_2_QN;
  (* src = "lattice_riscv.v:50722.6-50722.18" *)
  wire FD1P3BX_3_QN;
  (* src = "lattice_riscv.v:50725.6-50725.16" *)
  wire FD1P3BX_QN;
  wire GND_0_0_RED_VOTER_wire;
  (* src = "lattice_riscv.v:50721.6-50721.11" *)
  wire GND_0;
  (* src = "lattice_riscv.v:50721.6-50721.11" *)
  wire GND_0;
  (* src = "lattice_riscv.v:50721.6-50721.11" *)
  wire GND_0;
  (* src = "lattice_riscv.v:50630.6-50630.14" *)
  wire HFCLKCFG;
  (* src = "lattice_riscv.v:50631.6-50631.14" *)
  wire HFSDCOUT;
  (* src = "lattice_riscv.v:50632.6-50632.14" *)
  wire INTFBKOP;
  (* src = "lattice_riscv.v:50633.6-50633.14" *)
  wire INTFBKOS;
  (* src = "lattice_riscv.v:50634.6-50634.15" *)
  wire INTFBKOS2;
  (* src = "lattice_riscv.v:50635.6-50635.15" *)
  wire INTFBKOS3;
  (* src = "lattice_riscv.v:50636.6-50636.15" *)
  wire INTFBKOS4;
  (* src = "lattice_riscv.v:50637.6-50637.15" *)
  wire INTFBKOS5;
  (* src = "lattice_riscv.v:50644.6-50644.13" *)
  wire INTLOCK;
  (* src = "lattice_riscv.v:50645.6-50645.13" *)
  wire LEGRDYN;
  (* src = "lattice_riscv.v:50629.6-50629.14" *)
  wire LFCLKOUT;
  (* src = "lattice_riscv.v:50485.12-50485.21" *)
  wire [7:0] LMMIRDATA;
  (* src = "lattice_riscv.v:50638.6-50638.20" *)
  wire LMMIRDATAVALID;
  (* src = "lattice_riscv.v:50639.6-50639.15" *)
  wire LMMIREADY;
  (* src = "lattice_riscv.v:51254.6-51254.9" *)
  wire NC0;
  (* src = "lattice_riscv.v:50741.6-50741.11" *)
  wire N_100_TMR_0;
  (* src = "lattice_riscv.v:50741.6-50741.11" *)
  wire N_100_TMR_1;
  (* src = "lattice_riscv.v:50741.6-50741.11" *)
  wire N_100_TMR_2;
  wire N_103_0_RED_VOTER_wire;
  (* src = "lattice_riscv.v:50732.6-50732.11" *)
  wire N_103_TMR_0;
  (* src = "lattice_riscv.v:50732.6-50732.11" *)
  wire N_103_TMR_1;
  (* src = "lattice_riscv.v:50732.6-50732.11" *)
  wire N_103_TMR_2;
  (* src = "lattice_riscv.v:50739.6-50739.11" *)
  wire N_110_TMR_0;
  (* src = "lattice_riscv.v:50739.6-50739.11" *)
  wire N_110_TMR_1;
  (* src = "lattice_riscv.v:50739.6-50739.11" *)
  wire N_110_TMR_2;
  wire N_1209_i_0_RED_VOTER_wire;
  (* src = "lattice_riscv.v:51105.6-51105.14" *)
  wire N_1209_i_TMR_0;
  (* src = "lattice_riscv.v:51105.6-51105.14" *)
  wire N_1209_i_TMR_1;
  (* src = "lattice_riscv.v:51105.6-51105.14" *)
  wire N_1209_i_TMR_2;
  (* src = "lattice_riscv.v:51095.6-51095.13" *)
  wire N_120_i_TMR_0;
  (* src = "lattice_riscv.v:51095.6-51095.13" *)
  wire N_120_i_TMR_1;
  (* src = "lattice_riscv.v:51095.6-51095.13" *)
  wire N_120_i_TMR_2;
  (* src = "lattice_riscv.v:51100.6-51100.14" *)
  wire N_1210_i_TMR_0;
  (* src = "lattice_riscv.v:51100.6-51100.14" *)
  wire N_1210_i_TMR_1;
  (* src = "lattice_riscv.v:51100.6-51100.14" *)
  wire N_1210_i_TMR_2;
  (* src = "lattice_riscv.v:51178.6-51178.19" *)
  wire N_1210_i_fast_TMR_0;
  (* src = "lattice_riscv.v:51178.6-51178.19" *)
  wire N_1210_i_fast_TMR_1;
  (* src = "lattice_riscv.v:51178.6-51178.19" *)
  wire N_1210_i_fast_TMR_2;
  (* src = "lattice_riscv.v:51180.6-51180.19" *)
  wire N_1210_i_rep1_TMR_0;
  (* src = "lattice_riscv.v:51180.6-51180.19" *)
  wire N_1210_i_rep1_TMR_1;
  (* src = "lattice_riscv.v:51180.6-51180.19" *)
  wire N_1210_i_rep1_TMR_2;
  (* src = "lattice_riscv.v:51182.6-51182.19" *)
  wire N_1210_i_rep2_TMR_0;
  (* src = "lattice_riscv.v:51182.6-51182.19" *)
  wire N_1210_i_rep2_TMR_1;
  (* src = "lattice_riscv.v:51182.6-51182.19" *)
  wire N_1210_i_rep2_TMR_2;
  (* src = "lattice_riscv.v:51097.6-51097.14" *)
  wire N_1218_i_TMR_0;
  (* src = "lattice_riscv.v:51097.6-51097.14" *)
  wire N_1218_i_TMR_1;
  (* src = "lattice_riscv.v:51097.6-51097.14" *)
  wire N_1218_i_TMR_2;
  (* src = "lattice_riscv.v:51094.6-51094.14" *)
  wire N_1219_i_TMR_0;
  (* src = "lattice_riscv.v:51094.6-51094.14" *)
  wire N_1219_i_TMR_1;
  (* src = "lattice_riscv.v:51094.6-51094.14" *)
  wire N_1219_i_TMR_2;
  (* src = "lattice_riscv.v:51096.6-51096.13" *)
  wire N_121_i_TMR_0;
  (* src = "lattice_riscv.v:51096.6-51096.13" *)
  wire N_121_i_TMR_1;
  (* src = "lattice_riscv.v:51096.6-51096.13" *)
  wire N_121_i_TMR_2;
  (* src = "lattice_riscv.v:51098.6-51098.13" *)
  wire N_123_i_TMR_0;
  (* src = "lattice_riscv.v:51098.6-51098.13" *)
  wire N_123_i_TMR_1;
  (* src = "lattice_riscv.v:51098.6-51098.13" *)
  wire N_123_i_TMR_2;
  (* src = "lattice_riscv.v:51099.6-51099.13" *)
  wire N_124_i_TMR_0;
  (* src = "lattice_riscv.v:51099.6-51099.13" *)
  wire N_124_i_TMR_1;
  (* src = "lattice_riscv.v:51099.6-51099.13" *)
  wire N_124_i_TMR_2;
  (* src = "lattice_riscv.v:50860.6-50860.13" *)
  wire N_12821;
  (* src = "lattice_riscv.v:50861.6-50861.13" *)
  wire N_12822;
  (* src = "lattice_riscv.v:50862.6-50862.13" *)
  wire N_12823;
  (* src = "lattice_riscv.v:50863.6-50863.13" *)
  wire N_12824;
  (* src = "lattice_riscv.v:50864.6-50864.13" *)
  wire N_12825;
  (* src = "lattice_riscv.v:50865.6-50865.13" *)
  wire N_12826;
  (* src = "lattice_riscv.v:50866.6-50866.13" *)
  wire N_12827;
  (* src = "lattice_riscv.v:50867.6-50867.13" *)
  wire N_12828;
  (* src = "lattice_riscv.v:50868.6-50868.13" *)
  wire N_12829;
  (* src = "lattice_riscv.v:50869.6-50869.13" *)
  wire N_12830;
  (* src = "lattice_riscv.v:50870.6-50870.13" *)
  wire N_12831;
  (* src = "lattice_riscv.v:50871.6-50871.13" *)
  wire N_12832;
  (* src = "lattice_riscv.v:50872.6-50872.13" *)
  wire N_12833;
  (* src = "lattice_riscv.v:50873.6-50873.13" *)
  wire N_12834;
  (* src = "lattice_riscv.v:50874.6-50874.13" *)
  wire N_12835;
  (* src = "lattice_riscv.v:50875.6-50875.13" *)
  wire N_12836;
  (* src = "lattice_riscv.v:50876.6-50876.13" *)
  wire N_12837;
  (* src = "lattice_riscv.v:50877.6-50877.13" *)
  wire N_12838;
  (* src = "lattice_riscv.v:50878.6-50878.13" *)
  wire N_12839;
  (* src = "lattice_riscv.v:50879.6-50879.13" *)
  wire N_12840;
  (* src = "lattice_riscv.v:50880.6-50880.13" *)
  wire N_12841;
  (* src = "lattice_riscv.v:50881.6-50881.13" *)
  wire N_12842;
  (* src = "lattice_riscv.v:50882.6-50882.13" *)
  wire N_12843;
  (* src = "lattice_riscv.v:50883.6-50883.13" *)
  wire N_12844;
  (* src = "lattice_riscv.v:50884.6-50884.13" *)
  wire N_12845;
  (* src = "lattice_riscv.v:50885.6-50885.13" *)
  wire N_12846;
  (* src = "lattice_riscv.v:50886.6-50886.13" *)
  wire N_12847;
  (* src = "lattice_riscv.v:50887.6-50887.13" *)
  wire N_12848;
  (* src = "lattice_riscv.v:50888.6-50888.13" *)
  wire N_12849;
  (* src = "lattice_riscv.v:50889.6-50889.13" *)
  wire N_12850;
  (* src = "lattice_riscv.v:50890.6-50890.13" *)
  wire N_12851;
  (* src = "lattice_riscv.v:50891.6-50891.13" *)
  wire N_12852;
  (* src = "lattice_riscv.v:50892.6-50892.13" *)
  wire N_12853;
  (* src = "lattice_riscv.v:50893.6-50893.13" *)
  wire N_12854;
  (* src = "lattice_riscv.v:50894.6-50894.13" *)
  wire N_12855;
  (* src = "lattice_riscv.v:50895.6-50895.13" *)
  wire N_12856;
  (* src = "lattice_riscv.v:50896.6-50896.13" *)
  wire N_12857;
  (* src = "lattice_riscv.v:50897.6-50897.13" *)
  wire N_12858;
  (* src = "lattice_riscv.v:50898.6-50898.13" *)
  wire N_12859;
  (* src = "lattice_riscv.v:50899.6-50899.13" *)
  wire N_12860;
  (* src = "lattice_riscv.v:50900.6-50900.13" *)
  wire N_12861;
  (* src = "lattice_riscv.v:50901.6-50901.13" *)
  wire N_12862;
  (* src = "lattice_riscv.v:50902.6-50902.13" *)
  wire N_12863;
  (* src = "lattice_riscv.v:50903.6-50903.13" *)
  wire N_12864;
  (* src = "lattice_riscv.v:50904.6-50904.13" *)
  wire N_12865;
  (* src = "lattice_riscv.v:50905.6-50905.13" *)
  wire N_12866;
  (* src = "lattice_riscv.v:50906.6-50906.13" *)
  wire N_12867;
  (* src = "lattice_riscv.v:50907.6-50907.13" *)
  wire N_12868;
  (* src = "lattice_riscv.v:50908.6-50908.13" *)
  wire N_12869;
  (* src = "lattice_riscv.v:50909.6-50909.13" *)
  wire N_12870;
  (* src = "lattice_riscv.v:50910.6-50910.13" *)
  wire N_12871;
  (* src = "lattice_riscv.v:50911.6-50911.13" *)
  wire N_12872;
  (* src = "lattice_riscv.v:50912.6-50912.13" *)
  wire N_12873;
  (* src = "lattice_riscv.v:50913.6-50913.13" *)
  wire N_12874;
  (* src = "lattice_riscv.v:50914.6-50914.13" *)
  wire N_12875;
  (* src = "lattice_riscv.v:50915.6-50915.13" *)
  wire N_12876;
  (* src = "lattice_riscv.v:50916.6-50916.13" *)
  wire N_12877;
  (* src = "lattice_riscv.v:50917.6-50917.13" *)
  wire N_12878;
  (* src = "lattice_riscv.v:50918.6-50918.13" *)
  wire N_12879;
  (* src = "lattice_riscv.v:50919.6-50919.13" *)
  wire N_12880;
  (* src = "lattice_riscv.v:50920.6-50920.13" *)
  wire N_12881;
  (* src = "lattice_riscv.v:50921.6-50921.13" *)
  wire N_12882;
  (* src = "lattice_riscv.v:50922.6-50922.13" *)
  wire N_12883;
  (* src = "lattice_riscv.v:50923.6-50923.13" *)
  wire N_12884;
  (* src = "lattice_riscv.v:50924.6-50924.13" *)
  wire N_12885;
  (* src = "lattice_riscv.v:50925.6-50925.13" *)
  wire N_12886;
  (* src = "lattice_riscv.v:50926.6-50926.13" *)
  wire N_12887;
  (* src = "lattice_riscv.v:50927.6-50927.13" *)
  wire N_12888;
  (* src = "lattice_riscv.v:50928.6-50928.13" *)
  wire N_12889;
  (* src = "lattice_riscv.v:50929.6-50929.13" *)
  wire N_12890;
  (* src = "lattice_riscv.v:50930.6-50930.13" *)
  wire N_12891;
  (* src = "lattice_riscv.v:50931.6-50931.13" *)
  wire N_12892;
  (* src = "lattice_riscv.v:50932.6-50932.13" *)
  wire N_12893;
  (* src = "lattice_riscv.v:50933.6-50933.13" *)
  wire N_12894;
  (* src = "lattice_riscv.v:50934.6-50934.13" *)
  wire N_12895;
  (* src = "lattice_riscv.v:50935.6-50935.13" *)
  wire N_12896;
  (* src = "lattice_riscv.v:50936.6-50936.13" *)
  wire N_12897;
  (* src = "lattice_riscv.v:50937.6-50937.13" *)
  wire N_12898;
  (* src = "lattice_riscv.v:50938.6-50938.13" *)
  wire N_12899;
  (* src = "lattice_riscv.v:50939.6-50939.13" *)
  wire N_12900;
  (* src = "lattice_riscv.v:50940.6-50940.13" *)
  wire N_12901;
  (* src = "lattice_riscv.v:50941.6-50941.13" *)
  wire N_12902;
  (* src = "lattice_riscv.v:50942.6-50942.13" *)
  wire N_12903;
  (* src = "lattice_riscv.v:50943.6-50943.13" *)
  wire N_12904;
  (* src = "lattice_riscv.v:50944.6-50944.13" *)
  wire N_12905;
  (* src = "lattice_riscv.v:50945.6-50945.13" *)
  wire N_12906;
  (* src = "lattice_riscv.v:50946.6-50946.13" *)
  wire N_12907;
  (* src = "lattice_riscv.v:50947.6-50947.13" *)
  wire N_12908;
  (* src = "lattice_riscv.v:50948.6-50948.13" *)
  wire N_12909;
  (* src = "lattice_riscv.v:50949.6-50949.13" *)
  wire N_12910;
  (* src = "lattice_riscv.v:50950.6-50950.13" *)
  wire N_12911;
  (* src = "lattice_riscv.v:50951.6-50951.13" *)
  wire N_12912;
  (* src = "lattice_riscv.v:50952.6-50952.13" *)
  wire N_12913;
  (* src = "lattice_riscv.v:50953.6-50953.13" *)
  wire N_12914;
  (* src = "lattice_riscv.v:50954.6-50954.13" *)
  wire N_12915;
  (* src = "lattice_riscv.v:50955.6-50955.13" *)
  wire N_12916;
  (* src = "lattice_riscv.v:50956.6-50956.13" *)
  wire N_12917;
  (* src = "lattice_riscv.v:50957.6-50957.13" *)
  wire N_12918;
  (* src = "lattice_riscv.v:50958.6-50958.13" *)
  wire N_12919;
  (* src = "lattice_riscv.v:50959.6-50959.13" *)
  wire N_12920;
  (* src = "lattice_riscv.v:50960.6-50960.13" *)
  wire N_12921;
  (* src = "lattice_riscv.v:50961.6-50961.13" *)
  wire N_12922;
  (* src = "lattice_riscv.v:50962.6-50962.13" *)
  wire N_12923;
  (* src = "lattice_riscv.v:50963.6-50963.13" *)
  wire N_12924;
  (* src = "lattice_riscv.v:50964.6-50964.13" *)
  wire N_12925;
  (* src = "lattice_riscv.v:50965.6-50965.13" *)
  wire N_12926;
  (* src = "lattice_riscv.v:50966.6-50966.13" *)
  wire N_12927;
  (* src = "lattice_riscv.v:50967.6-50967.13" *)
  wire N_12928;
  (* src = "lattice_riscv.v:50968.6-50968.13" *)
  wire N_12929;
  (* src = "lattice_riscv.v:50969.6-50969.13" *)
  wire N_12930;
  (* src = "lattice_riscv.v:50970.6-50970.13" *)
  wire N_12931;
  (* src = "lattice_riscv.v:50971.6-50971.13" *)
  wire N_12932;
  (* src = "lattice_riscv.v:50972.6-50972.13" *)
  wire N_12933;
  (* src = "lattice_riscv.v:50973.6-50973.13" *)
  wire N_12934;
  (* src = "lattice_riscv.v:50974.6-50974.13" *)
  wire N_12935;
  (* src = "lattice_riscv.v:50975.6-50975.13" *)
  wire N_12936;
  (* src = "lattice_riscv.v:50976.6-50976.13" *)
  wire N_12937;
  (* src = "lattice_riscv.v:50977.6-50977.13" *)
  wire N_12938;
  (* src = "lattice_riscv.v:50978.6-50978.13" *)
  wire N_12939;
  (* src = "lattice_riscv.v:50979.6-50979.13" *)
  wire N_12940;
  (* src = "lattice_riscv.v:50980.6-50980.13" *)
  wire N_12941;
  (* src = "lattice_riscv.v:50981.6-50981.13" *)
  wire N_12942;
  (* src = "lattice_riscv.v:50982.6-50982.13" *)
  wire N_12943;
  (* src = "lattice_riscv.v:50983.6-50983.13" *)
  wire N_12944;
  (* src = "lattice_riscv.v:50984.6-50984.13" *)
  wire N_12945;
  (* src = "lattice_riscv.v:50985.6-50985.13" *)
  wire N_12946;
  (* src = "lattice_riscv.v:50740.6-50740.11" *)
  wire N_136_TMR_0;
  (* src = "lattice_riscv.v:50740.6-50740.11" *)
  wire N_136_TMR_1;
  (* src = "lattice_riscv.v:50740.6-50740.11" *)
  wire N_136_TMR_2;
  (* src = "lattice_riscv.v:51093.6-51093.13" *)
  wire N_137_i_TMR_0;
  (* src = "lattice_riscv.v:51093.6-51093.13" *)
  wire N_137_i_TMR_1;
  (* src = "lattice_riscv.v:51093.6-51093.13" *)
  wire N_137_i_TMR_2;
  (* src = "lattice_riscv.v:50742.6-50742.11" *)
  wire N_148_TMR_0;
  (* src = "lattice_riscv.v:50742.6-50742.11" *)
  wire N_148_TMR_1;
  (* src = "lattice_riscv.v:50742.6-50742.11" *)
  wire N_148_TMR_2;
  (* src = "lattice_riscv.v:51101.6-51101.13" *)
  wire N_152_i_TMR_0;
  (* src = "lattice_riscv.v:51101.6-51101.13" *)
  wire N_152_i_TMR_1;
  (* src = "lattice_riscv.v:51101.6-51101.13" *)
  wire N_152_i_TMR_2;
  (* src = "lattice_riscv.v:50743.6-50743.11" *)
  wire N_167_TMR_0;
  (* src = "lattice_riscv.v:50743.6-50743.11" *)
  wire N_167_TMR_1;
  (* src = "lattice_riscv.v:50743.6-50743.11" *)
  wire N_167_TMR_2;
  (* src = "lattice_riscv.v:50744.6-50744.11" *)
  wire N_175_TMR_0;
  (* src = "lattice_riscv.v:50744.6-50744.11" *)
  wire N_175_TMR_1;
  (* src = "lattice_riscv.v:50744.6-50744.11" *)
  wire N_175_TMR_2;
  (* src = "lattice_riscv.v:51245.6-51245.15" *)
  wire N_17815_0_TMR_0;
  (* src = "lattice_riscv.v:51245.6-51245.15" *)
  wire N_17815_0_TMR_1;
  (* src = "lattice_riscv.v:51245.6-51245.15" *)
  wire N_17815_0_TMR_2;
  (* src = "lattice_riscv.v:51244.6-51244.15" *)
  wire N_17817_0_TMR_0;
  (* src = "lattice_riscv.v:51244.6-51244.15" *)
  wire N_17817_0_TMR_1;
  (* src = "lattice_riscv.v:51244.6-51244.15" *)
  wire N_17817_0_TMR_2;
  (* src = "lattice_riscv.v:51243.6-51243.15" *)
  wire N_17819_0_TMR_0;
  (* src = "lattice_riscv.v:51243.6-51243.15" *)
  wire N_17819_0_TMR_1;
  (* src = "lattice_riscv.v:51243.6-51243.15" *)
  wire N_17819_0_TMR_2;
  (* src = "lattice_riscv.v:51242.6-51242.15" *)
  wire N_17821_0_TMR_0;
  (* src = "lattice_riscv.v:51242.6-51242.15" *)
  wire N_17821_0_TMR_1;
  (* src = "lattice_riscv.v:51242.6-51242.15" *)
  wire N_17821_0_TMR_2;
  (* src = "lattice_riscv.v:51241.6-51241.15" *)
  wire N_17823_0_TMR_0;
  (* src = "lattice_riscv.v:51241.6-51241.15" *)
  wire N_17823_0_TMR_1;
  (* src = "lattice_riscv.v:51241.6-51241.15" *)
  wire N_17823_0_TMR_2;
  (* src = "lattice_riscv.v:51240.6-51240.15" *)
  wire N_17825_0_TMR_0;
  (* src = "lattice_riscv.v:51240.6-51240.15" *)
  wire N_17825_0_TMR_1;
  (* src = "lattice_riscv.v:51240.6-51240.15" *)
  wire N_17825_0_TMR_2;
  (* src = "lattice_riscv.v:51239.6-51239.15" *)
  wire N_17827_0_TMR_0;
  (* src = "lattice_riscv.v:51239.6-51239.15" *)
  wire N_17827_0_TMR_1;
  (* src = "lattice_riscv.v:51239.6-51239.15" *)
  wire N_17827_0_TMR_2;
  (* src = "lattice_riscv.v:51238.6-51238.15" *)
  wire N_17829_0_TMR_0;
  (* src = "lattice_riscv.v:51238.6-51238.15" *)
  wire N_17829_0_TMR_1;
  (* src = "lattice_riscv.v:51238.6-51238.15" *)
  wire N_17829_0_TMR_2;
  (* src = "lattice_riscv.v:51237.6-51237.15" *)
  wire N_17831_0_TMR_0;
  (* src = "lattice_riscv.v:51237.6-51237.15" *)
  wire N_17831_0_TMR_1;
  (* src = "lattice_riscv.v:51237.6-51237.15" *)
  wire N_17831_0_TMR_2;
  (* src = "lattice_riscv.v:51236.6-51236.15" *)
  wire N_17833_0_TMR_0;
  (* src = "lattice_riscv.v:51236.6-51236.15" *)
  wire N_17833_0_TMR_1;
  (* src = "lattice_riscv.v:51236.6-51236.15" *)
  wire N_17833_0_TMR_2;
  (* src = "lattice_riscv.v:51235.6-51235.15" *)
  wire N_17835_0_TMR_0;
  (* src = "lattice_riscv.v:51235.6-51235.15" *)
  wire N_17835_0_TMR_1;
  (* src = "lattice_riscv.v:51235.6-51235.15" *)
  wire N_17835_0_TMR_2;
  (* src = "lattice_riscv.v:51234.6-51234.15" *)
  wire N_17837_0_TMR_0;
  (* src = "lattice_riscv.v:51234.6-51234.15" *)
  wire N_17837_0_TMR_1;
  (* src = "lattice_riscv.v:51234.6-51234.15" *)
  wire N_17837_0_TMR_2;
  (* src = "lattice_riscv.v:50737.6-50737.10" *)
  wire N_20_TMR_0;
  (* src = "lattice_riscv.v:50737.6-50737.10" *)
  wire N_20_TMR_1;
  (* src = "lattice_riscv.v:50737.6-50737.10" *)
  wire N_20_TMR_2;
  (* src = "lattice_riscv.v:51250.6-51250.13" *)
  wire N_22656;
  (* src = "lattice_riscv.v:51251.6-51251.13" *)
  wire N_22657_TMR_0;
  (* src = "lattice_riscv.v:51251.6-51251.13" *)
  wire N_22657_TMR_1;
  (* src = "lattice_riscv.v:51251.6-51251.13" *)
  wire N_22657_TMR_2;
  (* src = "lattice_riscv.v:51252.6-51252.13" *)
  wire N_22658;
  (* src = "lattice_riscv.v:51253.6-51253.13" *)
  wire N_22659_TMR_0;
  (* src = "lattice_riscv.v:51253.6-51253.13" *)
  wire N_22659_TMR_1;
  (* src = "lattice_riscv.v:51253.6-51253.13" *)
  wire N_22659_TMR_2;
  (* src = "lattice_riscv.v:50812.6-50812.11" *)
  wire N_403_TMR_0;
  (* src = "lattice_riscv.v:50812.6-50812.11" *)
  wire N_403_TMR_1;
  (* src = "lattice_riscv.v:50812.6-50812.11" *)
  wire N_403_TMR_2;
  (* src = "lattice_riscv.v:50813.6-50813.11" *)
  wire N_404_TMR_0;
  (* src = "lattice_riscv.v:50813.6-50813.11" *)
  wire N_404_TMR_1;
  (* src = "lattice_riscv.v:50813.6-50813.11" *)
  wire N_404_TMR_2;
  (* src = "lattice_riscv.v:50814.6-50814.11" *)
  wire N_405_TMR_0;
  (* src = "lattice_riscv.v:50814.6-50814.11" *)
  wire N_405_TMR_1;
  (* src = "lattice_riscv.v:50814.6-50814.11" *)
  wire N_405_TMR_2;
  (* src = "lattice_riscv.v:50815.6-50815.11" *)
  wire N_406_TMR_0;
  (* src = "lattice_riscv.v:50815.6-50815.11" *)
  wire N_406_TMR_1;
  (* src = "lattice_riscv.v:50815.6-50815.11" *)
  wire N_406_TMR_2;
  (* src = "lattice_riscv.v:50816.6-50816.11" *)
  wire N_407_TMR_0;
  (* src = "lattice_riscv.v:50816.6-50816.11" *)
  wire N_407_TMR_1;
  (* src = "lattice_riscv.v:50816.6-50816.11" *)
  wire N_407_TMR_2;
  (* src = "lattice_riscv.v:50817.6-50817.11" *)
  wire N_408_TMR_0;
  (* src = "lattice_riscv.v:50817.6-50817.11" *)
  wire N_408_TMR_1;
  (* src = "lattice_riscv.v:50817.6-50817.11" *)
  wire N_408_TMR_2;
  (* src = "lattice_riscv.v:50818.6-50818.11" *)
  wire N_409_TMR_0;
  (* src = "lattice_riscv.v:50818.6-50818.11" *)
  wire N_409_TMR_1;
  (* src = "lattice_riscv.v:50818.6-50818.11" *)
  wire N_409_TMR_2;
  (* src = "lattice_riscv.v:50819.6-50819.11" *)
  wire N_410_TMR_0;
  (* src = "lattice_riscv.v:50819.6-50819.11" *)
  wire N_410_TMR_1;
  (* src = "lattice_riscv.v:50819.6-50819.11" *)
  wire N_410_TMR_2;
  (* src = "lattice_riscv.v:50820.6-50820.11" *)
  wire N_411_TMR_0;
  (* src = "lattice_riscv.v:50820.6-50820.11" *)
  wire N_411_TMR_1;
  (* src = "lattice_riscv.v:50820.6-50820.11" *)
  wire N_411_TMR_2;
  (* src = "lattice_riscv.v:50821.6-50821.11" *)
  wire N_412_TMR_0;
  (* src = "lattice_riscv.v:50821.6-50821.11" *)
  wire N_412_TMR_1;
  (* src = "lattice_riscv.v:50821.6-50821.11" *)
  wire N_412_TMR_2;
  (* src = "lattice_riscv.v:50822.6-50822.11" *)
  wire N_413_TMR_0;
  (* src = "lattice_riscv.v:50822.6-50822.11" *)
  wire N_413_TMR_1;
  (* src = "lattice_riscv.v:50822.6-50822.11" *)
  wire N_413_TMR_2;
  (* src = "lattice_riscv.v:50823.6-50823.11" *)
  wire N_414_TMR_0;
  (* src = "lattice_riscv.v:50823.6-50823.11" *)
  wire N_414_TMR_1;
  (* src = "lattice_riscv.v:50823.6-50823.11" *)
  wire N_414_TMR_2;
  (* src = "lattice_riscv.v:50824.6-50824.11" *)
  wire N_415_TMR_0;
  (* src = "lattice_riscv.v:50824.6-50824.11" *)
  wire N_415_TMR_1;
  (* src = "lattice_riscv.v:50824.6-50824.11" *)
  wire N_415_TMR_2;
  (* src = "lattice_riscv.v:50825.6-50825.11" *)
  wire N_416_TMR_0;
  (* src = "lattice_riscv.v:50825.6-50825.11" *)
  wire N_416_TMR_1;
  (* src = "lattice_riscv.v:50825.6-50825.11" *)
  wire N_416_TMR_2;
  (* src = "lattice_riscv.v:50826.6-50826.11" *)
  wire N_417_TMR_0;
  (* src = "lattice_riscv.v:50826.6-50826.11" *)
  wire N_417_TMR_1;
  (* src = "lattice_riscv.v:50826.6-50826.11" *)
  wire N_417_TMR_2;
  (* src = "lattice_riscv.v:50828.6-50828.11" *)
  wire N_419_TMR_0;
  (* src = "lattice_riscv.v:50828.6-50828.11" *)
  wire N_419_TMR_1;
  (* src = "lattice_riscv.v:50828.6-50828.11" *)
  wire N_419_TMR_2;
  (* src = "lattice_riscv.v:50829.6-50829.11" *)
  wire N_420_TMR_0;
  (* src = "lattice_riscv.v:50829.6-50829.11" *)
  wire N_420_TMR_1;
  (* src = "lattice_riscv.v:50829.6-50829.11" *)
  wire N_420_TMR_2;
  (* src = "lattice_riscv.v:50832.6-50832.11" *)
  wire N_423_TMR_0;
  (* src = "lattice_riscv.v:50832.6-50832.11" *)
  wire N_423_TMR_1;
  (* src = "lattice_riscv.v:50832.6-50832.11" *)
  wire N_423_TMR_2;
  (* src = "lattice_riscv.v:50833.6-50833.11" *)
  wire N_424_TMR_0;
  (* src = "lattice_riscv.v:50833.6-50833.11" *)
  wire N_424_TMR_1;
  (* src = "lattice_riscv.v:50833.6-50833.11" *)
  wire N_424_TMR_2;
  (* src = "lattice_riscv.v:50834.6-50834.11" *)
  wire N_425_TMR_0;
  (* src = "lattice_riscv.v:50834.6-50834.11" *)
  wire N_425_TMR_1;
  (* src = "lattice_riscv.v:50834.6-50834.11" *)
  wire N_425_TMR_2;
  (* src = "lattice_riscv.v:50836.6-50836.11" *)
  wire N_427_TMR_0;
  (* src = "lattice_riscv.v:50836.6-50836.11" *)
  wire N_427_TMR_1;
  (* src = "lattice_riscv.v:50836.6-50836.11" *)
  wire N_427_TMR_2;
  (* src = "lattice_riscv.v:50837.6-50837.11" *)
  wire N_428_TMR_0;
  (* src = "lattice_riscv.v:50837.6-50837.11" *)
  wire N_428_TMR_1;
  (* src = "lattice_riscv.v:50837.6-50837.11" *)
  wire N_428_TMR_2;
  (* src = "lattice_riscv.v:50838.6-50838.11" *)
  wire N_429_TMR_0;
  (* src = "lattice_riscv.v:50838.6-50838.11" *)
  wire N_429_TMR_1;
  (* src = "lattice_riscv.v:50838.6-50838.11" *)
  wire N_429_TMR_2;
  (* src = "lattice_riscv.v:50839.6-50839.11" *)
  wire N_430_TMR_0;
  (* src = "lattice_riscv.v:50839.6-50839.11" *)
  wire N_430_TMR_1;
  (* src = "lattice_riscv.v:50839.6-50839.11" *)
  wire N_430_TMR_2;
  (* src = "lattice_riscv.v:50521.12-50521.17" *)
  wire N_443_TMR_0;
  (* src = "lattice_riscv.v:50521.12-50521.17" *)
  wire N_443_TMR_1;
  (* src = "lattice_riscv.v:50521.12-50521.17" *)
  wire N_443_TMR_2;
  (* src = "lattice_riscv.v:50769.6-50769.11" *)
  wire N_697_TMR_0;
  (* src = "lattice_riscv.v:50769.6-50769.11" *)
  wire N_697_TMR_1;
  (* src = "lattice_riscv.v:50769.6-50769.11" *)
  wire N_697_TMR_2;
  (* src = "lattice_riscv.v:50770.6-50770.11" *)
  wire N_698_TMR_0;
  (* src = "lattice_riscv.v:50770.6-50770.11" *)
  wire N_698_TMR_1;
  (* src = "lattice_riscv.v:50770.6-50770.11" *)
  wire N_698_TMR_2;
  (* src = "lattice_riscv.v:50771.6-50771.11" *)
  wire N_699_TMR_0;
  (* src = "lattice_riscv.v:50771.6-50771.11" *)
  wire N_699_TMR_1;
  (* src = "lattice_riscv.v:50771.6-50771.11" *)
  wire N_699_TMR_2;
  (* src = "lattice_riscv.v:50556.12-50556.17" *)
  wire N_792_TMR_0;
  (* src = "lattice_riscv.v:50556.12-50556.17" *)
  wire N_792_TMR_1;
  (* src = "lattice_riscv.v:50556.12-50556.17" *)
  wire N_792_TMR_2;
  (* src = "lattice_riscv.v:50738.6-50738.10" *)
  wire N_92_TMR_0;
  (* src = "lattice_riscv.v:50738.6-50738.10" *)
  wire N_92_TMR_1;
  (* src = "lattice_riscv.v:50738.6-50738.10" *)
  wire N_92_TMR_2;
  (* src = "lattice_riscv.v:50646.6-50646.11" *)
  wire PFDDN;
  (* src = "lattice_riscv.v:50647.6-50647.11" *)
  wire PFDUP;
  (* src = "lattice_riscv.v:50648.6-50648.14" *)
  wire REFMUXCK;
  (* src = "lattice_riscv.v:50649.6-50649.11" *)
  wire REGQA;
  (* src = "lattice_riscv.v:50650.6-50650.11" *)
  wire REGQB;
  (* src = "lattice_riscv.v:50651.6-50651.12" *)
  wire REGQB1;
  (* src = "lattice_riscv.v:50483.12-50483.28" *)
  wire [1:0] SP512K_1_ERRDECA;
  (* src = "lattice_riscv.v:50484.12-50484.28" *)
  wire [1:0] SP512K_1_ERRDECB;
  (* src = "lattice_riscv.v:50481.12-50481.26" *)
  wire [1:0] SP512K_ERRDECA;
  (* src = "lattice_riscv.v:50482.12-50482.26" *)
  wire [1:0] SP512K_ERRDECB;
  wire VCC_0_RED_VOTER_wire;
  (* src = "lattice_riscv.v:50628.6-50628.9" *)
  wire VCC_TMR_0;
  (* src = "lattice_riscv.v:50628.6-50628.9" *)
  wire VCC_TMR_1;
  (* src = "lattice_riscv.v:50628.6-50628.9" *)
  wire VCC_TMR_2;
  (* src = "lattice_riscv.v:51176.6-51176.100" *)
  wire \VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_0 ;
  (* src = "lattice_riscv.v:51176.6-51176.100" *)
  wire \VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_1 ;
  (* src = "lattice_riscv.v:51176.6-51176.100" *)
  wire \VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_2 ;
  (* src = "lattice_riscv.v:51088.6-51088.71" *)
  wire \VexRiscv.IBusCachedPlugin_cache.builder_slave_sel_r_r_0_a2_0_out_TMR_0 ;
  (* src = "lattice_riscv.v:51088.6-51088.71" *)
  wire \VexRiscv.IBusCachedPlugin_cache.builder_slave_sel_r_r_0_a2_0_out_TMR_1 ;
  (* src = "lattice_riscv.v:51088.6-51088.71" *)
  wire \VexRiscv.IBusCachedPlugin_cache.builder_slave_sel_r_r_0_a2_0_out_TMR_2 ;
  (* src = "lattice_riscv.v:50989.6-50989.69" *)
  wire \VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_0_0_TMR_0 ;
  (* src = "lattice_riscv.v:50989.6-50989.69" *)
  wire \VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_0_0_TMR_1 ;
  (* src = "lattice_riscv.v:50989.6-50989.69" *)
  wire \VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_0_0_TMR_2 ;
  (* src = "lattice_riscv.v:50539.13-50539.74" *)
  wire [31:1] \VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 ;
  (* src = "lattice_riscv.v:50539.13-50539.74" *)
  wire [31:1] \VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 ;
  (* src = "lattice_riscv.v:50539.13-50539.74" *)
  wire [31:1] \VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 ;
  (* src = "lattice_riscv.v:50538.13-50538.72" *)
  wire [31:1] \VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_0 ;
  (* src = "lattice_riscv.v:50538.13-50538.72" *)
  wire [31:1] \VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_1 ;
  (* src = "lattice_riscv.v:50538.13-50538.72" *)
  wire [31:1] \VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_2 ;
  (* src = "lattice_riscv.v:51144.6-51144.69" *)
  wire \VexRiscv.builder_csr_bankarray_interface0_bank_bus_dat_r10_3_0_TMR_0 ;
  (* src = "lattice_riscv.v:51144.6-51144.69" *)
  wire \VexRiscv.builder_csr_bankarray_interface0_bank_bus_dat_r10_3_0_TMR_1 ;
  (* src = "lattice_riscv.v:51144.6-51144.69" *)
  wire \VexRiscv.builder_csr_bankarray_interface0_bank_bus_dat_r10_3_0_TMR_2 ;
  (* src = "lattice_riscv.v:51087.6-51087.66" *)
  wire \VexRiscv.builder_csr_bankarray_interface0_bank_bus_dat_r8_0_TMR_0 ;
  (* src = "lattice_riscv.v:51087.6-51087.66" *)
  wire \VexRiscv.builder_csr_bankarray_interface0_bank_bus_dat_r8_0_TMR_1 ;
  (* src = "lattice_riscv.v:51087.6-51087.66" *)
  wire \VexRiscv.builder_csr_bankarray_interface0_bank_bus_dat_r8_0_TMR_2 ;
  (* src = "lattice_riscv.v:51143.6-51143.29" *)
  wire \VexRiscv.main_m1_e_0_1_TMR_0 ;
  (* src = "lattice_riscv.v:51143.6-51143.29" *)
  wire \VexRiscv.main_m1_e_0_1_TMR_1 ;
  (* src = "lattice_riscv.v:51143.6-51143.29" *)
  wire \VexRiscv.main_m1_e_0_1_TMR_2 ;
  wire builder_array_muxed0_0_RED_VOTER_wire;
  wire builder_array_muxed0_10_RED_VOTER_wire;
  wire builder_array_muxed0_11_RED_VOTER_wire;
  wire builder_array_muxed0_12_RED_VOTER_wire;
  wire builder_array_muxed0_13_RED_VOTER_wire;
  wire builder_array_muxed0_1_RED_VOTER_wire;
  wire builder_array_muxed0_2_RED_VOTER_wire;
  wire builder_array_muxed0_4_RED_VOTER_wire;
  wire builder_array_muxed0_5_RED_VOTER_wire;
  wire builder_array_muxed0_6_RED_VOTER_wire;
  wire builder_array_muxed0_7_RED_VOTER_wire;
  wire builder_array_muxed0_8_RED_VOTER_wire;
  wire builder_array_muxed0_9_RED_VOTER_wire;
  (* src = "lattice_riscv.v:50532.13-50532.33" *)
  wire [13:0] builder_array_muxed0_TMR_0;
  (* src = "lattice_riscv.v:50532.13-50532.33" *)
  wire [13:0] builder_array_muxed0_TMR_1;
  (* src = "lattice_riscv.v:50532.13-50532.33" *)
  wire [13:0] builder_array_muxed0_TMR_2;
  wire builder_array_muxed1_0_RED_VOTER_wire;
  wire builder_array_muxed1_10_RED_VOTER_wire;
  wire builder_array_muxed1_11_RED_VOTER_wire;
  wire builder_array_muxed1_12_RED_VOTER_wire;
  wire builder_array_muxed1_13_RED_VOTER_wire;
  wire builder_array_muxed1_14_RED_VOTER_wire;
  wire builder_array_muxed1_15_RED_VOTER_wire;
  wire builder_array_muxed1_16_RED_VOTER_wire;
  wire builder_array_muxed1_17_RED_VOTER_wire;
  wire builder_array_muxed1_18_RED_VOTER_wire;
  wire builder_array_muxed1_19_RED_VOTER_wire;
  wire builder_array_muxed1_1_RED_VOTER_wire;
  wire builder_array_muxed1_20_RED_VOTER_wire;
  wire builder_array_muxed1_21_RED_VOTER_wire;
  wire builder_array_muxed1_22_RED_VOTER_wire;
  wire builder_array_muxed1_23_RED_VOTER_wire;
  wire builder_array_muxed1_24_RED_VOTER_wire;
  wire builder_array_muxed1_25_RED_VOTER_wire;
  wire builder_array_muxed1_26_RED_VOTER_wire;
  wire builder_array_muxed1_27_RED_VOTER_wire;
  wire builder_array_muxed1_28_RED_VOTER_wire;
  wire builder_array_muxed1_29_RED_VOTER_wire;
  wire builder_array_muxed1_2_RED_VOTER_wire;
  wire builder_array_muxed1_30_RED_VOTER_wire;
  wire builder_array_muxed1_31_RED_VOTER_wire;
  wire builder_array_muxed1_3_RED_VOTER_wire;
  wire builder_array_muxed1_4_RED_VOTER_wire;
  wire builder_array_muxed1_5_RED_VOTER_wire;
  wire builder_array_muxed1_6_RED_VOTER_wire;
  wire builder_array_muxed1_7_RED_VOTER_wire;
  wire builder_array_muxed1_8_RED_VOTER_wire;
  wire builder_array_muxed1_9_RED_VOTER_wire;
  (* src = "lattice_riscv.v:50486.13-50486.33" *)
  wire [31:0] builder_array_muxed1_TMR_0;
  (* src = "lattice_riscv.v:50486.13-50486.33" *)
  wire [31:0] builder_array_muxed1_TMR_1;
  (* src = "lattice_riscv.v:50486.13-50486.33" *)
  wire [31:0] builder_array_muxed1_TMR_2;
  wire builder_array_muxed2_i_0_RED_VOTER_wire;
  wire builder_array_muxed2_i_1_RED_VOTER_wire;
  wire builder_array_muxed2_i_2_RED_VOTER_wire;
  wire builder_array_muxed2_i_3_RED_VOTER_wire;
  (* src = "lattice_riscv.v:50563.12-50563.34" *)
  wire [3:0] builder_array_muxed2_i_TMR_0;
  (* src = "lattice_riscv.v:50563.12-50563.34" *)
  wire [3:0] builder_array_muxed2_i_TMR_1;
  (* src = "lattice_riscv.v:50563.12-50563.34" *)
  wire [3:0] builder_array_muxed2_i_TMR_2;
  (* src = "lattice_riscv.v:50520.12-50520.31" *)
  wire [5:0] builder_basesoc_adr_TMR_0;
  (* src = "lattice_riscv.v:50520.12-50520.31" *)
  wire [5:0] builder_basesoc_adr_TMR_1;
  (* src = "lattice_riscv.v:50520.12-50520.31" *)
  wire [5:0] builder_basesoc_adr_TMR_2;
  (* src = "lattice_riscv.v:50657.6-50657.27" *)
  wire builder_basesoc_clkfb;
  (* src = "lattice_riscv.v:50701.6-50701.43" *)
  wire builder_basesoc_next_state_1_sqmuxa_1_TMR_0;
  (* src = "lattice_riscv.v:50701.6-50701.43" *)
  wire builder_basesoc_next_state_1_sqmuxa_1_TMR_1;
  (* src = "lattice_riscv.v:50701.6-50701.43" *)
  wire builder_basesoc_next_state_1_sqmuxa_1_TMR_2;
  (* src = "lattice_riscv.v:51202.6-51202.41" *)
  wire builder_basesoc_rs232phyrx_state_QN;
  (* src = "lattice_riscv.v:50667.6-50667.38" *)
  wire builder_basesoc_rs232phyrx_state_TMR_0;
  (* src = "lattice_riscv.v:50667.6-50667.38" *)
  wire builder_basesoc_rs232phyrx_state_TMR_1;
  (* src = "lattice_riscv.v:50667.6-50667.38" *)
  wire builder_basesoc_rs232phyrx_state_TMR_2;
  (* src = "lattice_riscv.v:51248.6-51248.40" *)
  wire builder_basesoc_rs232phyrx_state_i_TMR_0;
  (* src = "lattice_riscv.v:51248.6-51248.40" *)
  wire builder_basesoc_rs232phyrx_state_i_TMR_1;
  (* src = "lattice_riscv.v:51248.6-51248.40" *)
  wire builder_basesoc_rs232phyrx_state_i_TMR_2;
  (* src = "lattice_riscv.v:51203.6-51203.41" *)
  wire builder_basesoc_rs232phytx_state_QN;
  (* src = "lattice_riscv.v:50666.6-50666.38" *)
  wire builder_basesoc_rs232phytx_state_TMR_0;
  (* src = "lattice_riscv.v:50666.6-50666.38" *)
  wire builder_basesoc_rs232phytx_state_TMR_1;
  (* src = "lattice_riscv.v:50666.6-50666.38" *)
  wire builder_basesoc_rs232phytx_state_TMR_2;
  (* src = "lattice_riscv.v:51249.6-51249.40" *)
  wire builder_basesoc_rs232phytx_state_i_TMR_0;
  (* src = "lattice_riscv.v:51249.6-51249.40" *)
  wire builder_basesoc_rs232phytx_state_i_TMR_1;
  (* src = "lattice_riscv.v:51249.6-51249.40" *)
  wire builder_basesoc_rs232phytx_state_i_TMR_2;
  (* src = "lattice_riscv.v:51204.6-51204.30" *)
  wire builder_basesoc_state_QN;
  (* src = "lattice_riscv.v:50670.6-50670.27" *)
  wire builder_basesoc_state_TMR_0;
  (* src = "lattice_riscv.v:50670.6-50670.27" *)
  wire builder_basesoc_state_TMR_1;
  (* src = "lattice_riscv.v:50670.6-50670.27" *)
  wire builder_basesoc_state_TMR_2;
  (* src = "lattice_riscv.v:50584.12-50584.34" *)
  wire [5:0] builder_count_0_mod_QN;
  (* src = "lattice_riscv.v:50548.12-50548.35" *)
  wire [5:0] builder_count_0_mod_RNO_TMR_0;
  (* src = "lattice_riscv.v:50548.12-50548.35" *)
  wire [5:0] builder_count_0_mod_RNO_TMR_1;
  (* src = "lattice_riscv.v:50548.12-50548.35" *)
  wire [5:0] builder_count_0_mod_RNO_TMR_2;
  (* src = "lattice_riscv.v:50557.13-50557.30" *)
  wire [19:6] builder_count_1_2_TMR_0;
  (* src = "lattice_riscv.v:50557.13-50557.30" *)
  wire [19:6] builder_count_1_2_TMR_1;
  (* src = "lattice_riscv.v:50557.13-50557.30" *)
  wire [19:6] builder_count_1_2_TMR_2;
  (* src = "lattice_riscv.v:50990.6-50990.21" *)
  wire builder_count_1_TMR_0;
  (* src = "lattice_riscv.v:50990.6-50990.21" *)
  wire builder_count_1_TMR_1;
  (* src = "lattice_riscv.v:50990.6-50990.21" *)
  wire builder_count_1_TMR_2;
  (* src = "lattice_riscv.v:51157.6-51157.32" *)
  wire builder_count_1_cry_0_0_S0_TMR_0;
  (* src = "lattice_riscv.v:51157.6-51157.32" *)
  wire builder_count_1_cry_0_0_S0_TMR_1;
  (* src = "lattice_riscv.v:51157.6-51157.32" *)
  wire builder_count_1_cry_0_0_S0_TMR_2;
  (* src = "lattice_riscv.v:51149.6-51149.32" *)
  wire builder_count_1_cry_0_0_S1_TMR_0;
  (* src = "lattice_riscv.v:51149.6-51149.32" *)
  wire builder_count_1_cry_0_0_S1_TMR_1;
  (* src = "lattice_riscv.v:51149.6-51149.32" *)
  wire builder_count_1_cry_0_0_S1_TMR_2;
  (* src = "lattice_riscv.v:51051.6-51051.27" *)
  wire builder_count_1_cry_0_TMR_0;
  (* src = "lattice_riscv.v:51051.6-51051.27" *)
  wire builder_count_1_cry_0_TMR_1;
  (* src = "lattice_riscv.v:51051.6-51051.27" *)
  wire builder_count_1_cry_0_TMR_2;
  (* src = "lattice_riscv.v:51056.6-51056.28" *)
  wire builder_count_1_cry_10_TMR_0;
  (* src = "lattice_riscv.v:51056.6-51056.28" *)
  wire builder_count_1_cry_10_TMR_1;
  (* src = "lattice_riscv.v:51056.6-51056.28" *)
  wire builder_count_1_cry_10_TMR_2;
  (* src = "lattice_riscv.v:50776.6-50776.33" *)
  wire builder_count_1_cry_11_0_S0_TMR_0;
  (* src = "lattice_riscv.v:50776.6-50776.33" *)
  wire builder_count_1_cry_11_0_S0_TMR_1;
  (* src = "lattice_riscv.v:50776.6-50776.33" *)
  wire builder_count_1_cry_11_0_S0_TMR_2;
  (* src = "lattice_riscv.v:50777.6-50777.33" *)
  wire builder_count_1_cry_11_0_S1_TMR_0;
  (* src = "lattice_riscv.v:50777.6-50777.33" *)
  wire builder_count_1_cry_11_0_S1_TMR_1;
  (* src = "lattice_riscv.v:50777.6-50777.33" *)
  wire builder_count_1_cry_11_0_S1_TMR_2;
  (* src = "lattice_riscv.v:51057.6-51057.28" *)
  wire builder_count_1_cry_12_TMR_0;
  (* src = "lattice_riscv.v:51057.6-51057.28" *)
  wire builder_count_1_cry_12_TMR_1;
  (* src = "lattice_riscv.v:51057.6-51057.28" *)
  wire builder_count_1_cry_12_TMR_2;
  (* src = "lattice_riscv.v:50778.6-50778.33" *)
  wire builder_count_1_cry_13_0_S0_TMR_0;
  (* src = "lattice_riscv.v:50778.6-50778.33" *)
  wire builder_count_1_cry_13_0_S0_TMR_1;
  (* src = "lattice_riscv.v:50778.6-50778.33" *)
  wire builder_count_1_cry_13_0_S0_TMR_2;
  (* src = "lattice_riscv.v:51058.6-51058.28" *)
  wire builder_count_1_cry_14_TMR_0;
  (* src = "lattice_riscv.v:51058.6-51058.28" *)
  wire builder_count_1_cry_14_TMR_1;
  (* src = "lattice_riscv.v:51058.6-51058.28" *)
  wire builder_count_1_cry_14_TMR_2;
  (* src = "lattice_riscv.v:50779.6-50779.33" *)
  wire builder_count_1_cry_15_0_S0_TMR_0;
  (* src = "lattice_riscv.v:50779.6-50779.33" *)
  wire builder_count_1_cry_15_0_S0_TMR_1;
  (* src = "lattice_riscv.v:50779.6-50779.33" *)
  wire builder_count_1_cry_15_0_S0_TMR_2;
  (* src = "lattice_riscv.v:51059.6-51059.28" *)
  wire builder_count_1_cry_16_TMR_0;
  (* src = "lattice_riscv.v:51059.6-51059.28" *)
  wire builder_count_1_cry_16_TMR_1;
  (* src = "lattice_riscv.v:51059.6-51059.28" *)
  wire builder_count_1_cry_16_TMR_2;
  (* src = "lattice_riscv.v:51060.6-51060.28" *)
  wire builder_count_1_cry_18_TMR_0;
  (* src = "lattice_riscv.v:51060.6-51060.28" *)
  wire builder_count_1_cry_18_TMR_1;
  (* src = "lattice_riscv.v:51060.6-51060.28" *)
  wire builder_count_1_cry_18_TMR_2;
  (* src = "lattice_riscv.v:50768.6-50768.32" *)
  wire builder_count_1_cry_1_0_S0_TMR_0;
  (* src = "lattice_riscv.v:50768.6-50768.32" *)
  wire builder_count_1_cry_1_0_S0_TMR_1;
  (* src = "lattice_riscv.v:50768.6-50768.32" *)
  wire builder_count_1_cry_1_0_S0_TMR_2;
  (* src = "lattice_riscv.v:51052.6-51052.27" *)
  wire builder_count_1_cry_2_TMR_0;
  (* src = "lattice_riscv.v:51052.6-51052.27" *)
  wire builder_count_1_cry_2_TMR_1;
  (* src = "lattice_riscv.v:51052.6-51052.27" *)
  wire builder_count_1_cry_2_TMR_2;
  (* src = "lattice_riscv.v:51053.6-51053.27" *)
  wire builder_count_1_cry_4_TMR_0;
  (* src = "lattice_riscv.v:51053.6-51053.27" *)
  wire builder_count_1_cry_4_TMR_1;
  (* src = "lattice_riscv.v:51053.6-51053.27" *)
  wire builder_count_1_cry_4_TMR_2;
  (* src = "lattice_riscv.v:50772.6-50772.32" *)
  wire builder_count_1_cry_5_0_S0_TMR_0;
  (* src = "lattice_riscv.v:50772.6-50772.32" *)
  wire builder_count_1_cry_5_0_S0_TMR_1;
  (* src = "lattice_riscv.v:50772.6-50772.32" *)
  wire builder_count_1_cry_5_0_S0_TMR_2;
  (* src = "lattice_riscv.v:51054.6-51054.27" *)
  wire builder_count_1_cry_6_TMR_0;
  (* src = "lattice_riscv.v:51054.6-51054.27" *)
  wire builder_count_1_cry_6_TMR_1;
  (* src = "lattice_riscv.v:51054.6-51054.27" *)
  wire builder_count_1_cry_6_TMR_2;
  (* src = "lattice_riscv.v:50773.6-50773.32" *)
  wire builder_count_1_cry_7_0_S0_TMR_0;
  (* src = "lattice_riscv.v:50773.6-50773.32" *)
  wire builder_count_1_cry_7_0_S0_TMR_1;
  (* src = "lattice_riscv.v:50773.6-50773.32" *)
  wire builder_count_1_cry_7_0_S0_TMR_2;
  (* src = "lattice_riscv.v:50774.6-50774.32" *)
  wire builder_count_1_cry_7_0_S1_TMR_0;
  (* src = "lattice_riscv.v:50774.6-50774.32" *)
  wire builder_count_1_cry_7_0_S1_TMR_1;
  (* src = "lattice_riscv.v:50774.6-50774.32" *)
  wire builder_count_1_cry_7_0_S1_TMR_2;
  (* src = "lattice_riscv.v:51055.6-51055.27" *)
  wire builder_count_1_cry_8_TMR_0;
  (* src = "lattice_riscv.v:51055.6-51055.27" *)
  wire builder_count_1_cry_8_TMR_1;
  (* src = "lattice_riscv.v:51055.6-51055.27" *)
  wire builder_count_1_cry_8_TMR_2;
  (* src = "lattice_riscv.v:50775.6-50775.32" *)
  wire builder_count_1_cry_9_0_S1_TMR_0;
  (* src = "lattice_riscv.v:50775.6-50775.32" *)
  wire builder_count_1_cry_9_0_S1_TMR_1;
  (* src = "lattice_riscv.v:50775.6-50775.32" *)
  wire builder_count_1_cry_9_0_S1_TMR_2;
  (* src = "lattice_riscv.v:51159.6-51159.33" *)
  wire builder_count_1_s_19_0_COUT_TMR_0;
  (* src = "lattice_riscv.v:51159.6-51159.33" *)
  wire builder_count_1_s_19_0_COUT_TMR_1;
  (* src = "lattice_riscv.v:51159.6-51159.33" *)
  wire builder_count_1_s_19_0_COUT_TMR_2;
  (* src = "lattice_riscv.v:51158.6-51158.31" *)
  wire builder_count_1_s_19_0_S1_TMR_0;
  (* src = "lattice_riscv.v:51158.6-51158.31" *)
  wire builder_count_1_s_19_0_S1_TMR_1;
  (* src = "lattice_riscv.v:51158.6-51158.31" *)
  wire builder_count_1_s_19_0_S1_TMR_2;
  (* src = "lattice_riscv.v:50583.13-50583.29" *)
  wire [19:6] builder_count_QN;
  (* src = "lattice_riscv.v:50585.12-50585.32" *)
  wire [4:2] builder_count_mod_QN;
  (* src = "lattice_riscv.v:50547.12-50547.33" *)
  wire [4:2] builder_count_mod_RNO_TMR_0;
  (* src = "lattice_riscv.v:50547.12-50547.33" *)
  wire [4:2] builder_count_mod_RNO_TMR_1;
  (* src = "lattice_riscv.v:50547.12-50547.33" *)
  wire [4:2] builder_count_mod_RNO_TMR_2;
  (* src = "lattice_riscv.v:50529.14-50529.29" *)
  wire [15:12] builder_count_r_TMR_0;
  (* src = "lattice_riscv.v:50529.14-50529.29" *)
  wire [15:12] builder_count_r_TMR_1;
  (* src = "lattice_riscv.v:50529.14-50529.29" *)
  wire [15:12] builder_count_r_TMR_2;
  (* src = "lattice_riscv.v:50702.6-50702.46" *)
  wire builder_csr_bankarray_csrbank0_reset0_re_TMR_0;
  (* src = "lattice_riscv.v:50702.6-50702.46" *)
  wire builder_csr_bankarray_csrbank0_reset0_re_TMR_1;
  (* src = "lattice_riscv.v:50702.6-50702.46" *)
  wire builder_csr_bankarray_csrbank0_reset0_re_TMR_2;
  (* src = "lattice_riscv.v:50703.6-50703.48" *)
  wire builder_csr_bankarray_csrbank0_scratch0_re_TMR_0;
  (* src = "lattice_riscv.v:50703.6-50703.48" *)
  wire builder_csr_bankarray_csrbank0_scratch0_re_TMR_1;
  (* src = "lattice_riscv.v:50703.6-50703.48" *)
  wire builder_csr_bankarray_csrbank0_scratch0_re_TMR_2;
  (* src = "lattice_riscv.v:50704.6-50704.44" *)
  wire builder_csr_bankarray_csrbank1_out0_re_TMR_0;
  (* src = "lattice_riscv.v:50704.6-50704.44" *)
  wire builder_csr_bankarray_csrbank1_out0_re_TMR_1;
  (* src = "lattice_riscv.v:50704.6-50704.44" *)
  wire builder_csr_bankarray_csrbank1_out0_re_TMR_2;
  (* src = "lattice_riscv.v:50706.6-50706.43" *)
  wire builder_csr_bankarray_csrbank2_en0_re_TMR_0;
  (* src = "lattice_riscv.v:50706.6-50706.43" *)
  wire builder_csr_bankarray_csrbank2_en0_re_TMR_1;
  (* src = "lattice_riscv.v:50706.6-50706.43" *)
  wire builder_csr_bankarray_csrbank2_en0_re_TMR_2;
  (* src = "lattice_riscv.v:50709.6-50709.50" *)
  wire builder_csr_bankarray_csrbank2_ev_enable0_re_TMR_0;
  (* src = "lattice_riscv.v:50709.6-50709.50" *)
  wire builder_csr_bankarray_csrbank2_ev_enable0_re_TMR_1;
  (* src = "lattice_riscv.v:50709.6-50709.50" *)
  wire builder_csr_bankarray_csrbank2_ev_enable0_re_TMR_2;
  (* src = "lattice_riscv.v:50708.6-50708.50" *)
  wire builder_csr_bankarray_csrbank2_ev_pending_re_TMR_0;
  (* src = "lattice_riscv.v:50708.6-50708.50" *)
  wire builder_csr_bankarray_csrbank2_ev_pending_re_TMR_1;
  (* src = "lattice_riscv.v:50708.6-50708.50" *)
  wire builder_csr_bankarray_csrbank2_ev_pending_re_TMR_2;
  (* src = "lattice_riscv.v:50705.6-50705.47" *)
  wire builder_csr_bankarray_csrbank2_reload0_re_TMR_0;
  (* src = "lattice_riscv.v:50705.6-50705.47" *)
  wire builder_csr_bankarray_csrbank2_reload0_re_TMR_1;
  (* src = "lattice_riscv.v:50705.6-50705.47" *)
  wire builder_csr_bankarray_csrbank2_reload0_re_TMR_2;
  (* src = "lattice_riscv.v:50707.6-50707.53" *)
  wire builder_csr_bankarray_csrbank2_update_value0_re_TMR_0;
  (* src = "lattice_riscv.v:50707.6-50707.53" *)
  wire builder_csr_bankarray_csrbank2_update_value0_re_TMR_1;
  (* src = "lattice_riscv.v:50707.6-50707.53" *)
  wire builder_csr_bankarray_csrbank2_update_value0_re_TMR_2;
  (* src = "lattice_riscv.v:50711.6-50711.50" *)
  wire builder_csr_bankarray_csrbank3_ev_enable0_re_TMR_0;
  (* src = "lattice_riscv.v:50711.6-50711.50" *)
  wire builder_csr_bankarray_csrbank3_ev_enable0_re_TMR_1;
  (* src = "lattice_riscv.v:50711.6-50711.50" *)
  wire builder_csr_bankarray_csrbank3_ev_enable0_re_TMR_2;
  (* src = "lattice_riscv.v:50710.6-50710.50" *)
  wire builder_csr_bankarray_csrbank3_ev_pending_re_TMR_0;
  (* src = "lattice_riscv.v:50710.6-50710.50" *)
  wire builder_csr_bankarray_csrbank3_ev_pending_re_TMR_1;
  (* src = "lattice_riscv.v:50710.6-50710.50" *)
  wire builder_csr_bankarray_csrbank3_ev_pending_re_TMR_2;
  (* src = "lattice_riscv.v:50734.6-50734.40" *)
  wire builder_csr_bankarray_csrbank3_sel_TMR_0;
  (* src = "lattice_riscv.v:50734.6-50734.40" *)
  wire builder_csr_bankarray_csrbank3_sel_TMR_1;
  (* src = "lattice_riscv.v:50734.6-50734.40" *)
  wire builder_csr_bankarray_csrbank3_sel_TMR_2;
  (* src = "lattice_riscv.v:51111.6-51111.46" *)
  wire \builder_csr_bankarray_dat_r_7_1_.N_13_i_TMR_0 ;
  (* src = "lattice_riscv.v:51111.6-51111.46" *)
  wire \builder_csr_bankarray_dat_r_7_1_.N_13_i_TMR_1 ;
  (* src = "lattice_riscv.v:51111.6-51111.46" *)
  wire \builder_csr_bankarray_dat_r_7_1_.N_13_i_TMR_2 ;
  (* src = "lattice_riscv.v:51114.6-51114.48" *)
  wire \builder_csr_bankarray_dat_r_7_1_.i2_mux_0_TMR_0 ;
  (* src = "lattice_riscv.v:51114.6-51114.48" *)
  wire \builder_csr_bankarray_dat_r_7_1_.i2_mux_0_TMR_1 ;
  (* src = "lattice_riscv.v:51114.6-51114.48" *)
  wire \builder_csr_bankarray_dat_r_7_1_.i2_mux_0_TMR_2 ;
  (* src = "lattice_riscv.v:51128.6-51128.48" *)
  wire \builder_csr_bankarray_dat_r_7_1_.i3_mux_3_TMR_0 ;
  (* src = "lattice_riscv.v:51128.6-51128.48" *)
  wire \builder_csr_bankarray_dat_r_7_1_.i3_mux_3_TMR_1 ;
  (* src = "lattice_riscv.v:51128.6-51128.48" *)
  wire \builder_csr_bankarray_dat_r_7_1_.i3_mux_3_TMR_2 ;
  (* src = "lattice_riscv.v:51129.6-51129.46" *)
  wire \builder_csr_bankarray_dat_r_7_1_.i4_mux_TMR_0 ;
  (* src = "lattice_riscv.v:51129.6-51129.46" *)
  wire \builder_csr_bankarray_dat_r_7_1_.i4_mux_TMR_1 ;
  (* src = "lattice_riscv.v:51129.6-51129.46" *)
  wire \builder_csr_bankarray_dat_r_7_1_.i4_mux_TMR_2 ;
  (* src = "lattice_riscv.v:51175.6-51175.48" *)
  wire \builder_csr_bankarray_dat_r_7_1_.m35_am_1_TMR_0 ;
  (* src = "lattice_riscv.v:51175.6-51175.48" *)
  wire \builder_csr_bankarray_dat_r_7_1_.m35_am_1_TMR_1 ;
  (* src = "lattice_riscv.v:51175.6-51175.48" *)
  wire \builder_csr_bankarray_dat_r_7_1_.m35_am_1_TMR_2 ;
  (* src = "lattice_riscv.v:50581.12-50581.39" *)
  wire [7:1] builder_csr_bankarray_dat_r_TMR_0;
  (* src = "lattice_riscv.v:50581.12-50581.39" *)
  wire [7:1] builder_csr_bankarray_dat_r_TMR_1;
  (* src = "lattice_riscv.v:50581.12-50581.39" *)
  wire [7:1] builder_csr_bankarray_dat_r_TMR_2;
  (* src = "lattice_riscv.v:51090.6-51090.65" *)
  wire builder_csr_bankarray_interface0_bank_bus_dat_r8_6_RNIG6FO8_TMR_0;
  (* src = "lattice_riscv.v:51090.6-51090.65" *)
  wire builder_csr_bankarray_interface0_bank_bus_dat_r8_6_RNIG6FO8_TMR_1;
  (* src = "lattice_riscv.v:51090.6-51090.65" *)
  wire builder_csr_bankarray_interface0_bank_bus_dat_r8_6_RNIG6FO8_TMR_2;
  (* src = "lattice_riscv.v:50531.13-50531.62" *)
  wire [31:0] builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_0;
  (* src = "lattice_riscv.v:50531.13-50531.62" *)
  wire [31:0] builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_1;
  (* src = "lattice_riscv.v:50531.13-50531.62" *)
  wire [31:0] builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_2;
  (* src = "lattice_riscv.v:50586.13-50586.63" *)
  wire [31:0] builder_csr_bankarray_interface0_bank_bus_dat_r_QN;
  (* src = "lattice_riscv.v:50499.13-50499.60" *)
  wire [31:0] builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_0;
  (* src = "lattice_riscv.v:50499.13-50499.60" *)
  wire [31:0] builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_1;
  (* src = "lattice_riscv.v:50499.13-50499.60" *)
  wire [31:0] builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_2;
  (* src = "lattice_riscv.v:51104.6-51104.64" *)
  wire builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_0;
  (* src = "lattice_riscv.v:51104.6-51104.64" *)
  wire builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_1;
  (* src = "lattice_riscv.v:51104.6-51104.64" *)
  wire builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_2;
  (* src = "lattice_riscv.v:50587.13-50587.63" *)
  wire [13:0] builder_csr_bankarray_interface1_bank_bus_dat_r_QN;
  (* src = "lattice_riscv.v:50500.13-50500.60" *)
  wire [13:0] builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_0;
  (* src = "lattice_riscv.v:50500.13-50500.60" *)
  wire [13:0] builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_1;
  (* src = "lattice_riscv.v:50500.13-50500.60" *)
  wire [13:0] builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_2;
  (* src = "lattice_riscv.v:50526.13-50526.63" *)
  wire [31:0] builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_0;
  (* src = "lattice_riscv.v:50526.13-50526.63" *)
  wire [31:0] builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_1;
  (* src = "lattice_riscv.v:50526.13-50526.63" *)
  wire [31:0] builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_2;
  (* src = "lattice_riscv.v:50588.13-50588.63" *)
  wire [31:0] builder_csr_bankarray_interface2_bank_bus_dat_r_QN;
  (* src = "lattice_riscv.v:50509.13-50509.60" *)
  wire [31:0] builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_0;
  (* src = "lattice_riscv.v:50509.13-50509.60" *)
  wire [31:0] builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_1;
  (* src = "lattice_riscv.v:50509.13-50509.60" *)
  wire [31:0] builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_2;
  (* src = "lattice_riscv.v:50733.6-50733.62" *)
  wire builder_csr_bankarray_interface3_bank_bus_dat_r_0_sqmuxa_TMR_0;
  (* src = "lattice_riscv.v:50733.6-50733.62" *)
  wire builder_csr_bankarray_interface3_bank_bus_dat_r_0_sqmuxa_TMR_1;
  (* src = "lattice_riscv.v:50733.6-50733.62" *)
  wire builder_csr_bankarray_interface3_bank_bus_dat_r_0_sqmuxa_TMR_2;
  (* src = "lattice_riscv.v:51102.6-51102.64" *)
  wire builder_csr_bankarray_interface3_bank_bus_dat_r_0_sqmuxa_i_TMR_0;
  (* src = "lattice_riscv.v:51102.6-51102.64" *)
  wire builder_csr_bankarray_interface3_bank_bus_dat_r_0_sqmuxa_i_TMR_1;
  (* src = "lattice_riscv.v:51102.6-51102.64" *)
  wire builder_csr_bankarray_interface3_bank_bus_dat_r_0_sqmuxa_i_TMR_2;
  (* src = "lattice_riscv.v:50527.12-50527.62" *)
  wire [1:0] builder_csr_bankarray_interface3_bank_bus_dat_r_11_TMR_0;
  (* src = "lattice_riscv.v:50527.12-50527.62" *)
  wire [1:0] builder_csr_bankarray_interface3_bank_bus_dat_r_11_TMR_1;
  (* src = "lattice_riscv.v:50527.12-50527.62" *)
  wire [1:0] builder_csr_bankarray_interface3_bank_bus_dat_r_11_TMR_2;
  (* src = "lattice_riscv.v:50589.12-50589.62" *)
  wire [7:0] builder_csr_bankarray_interface3_bank_bus_dat_r_QN;
  (* src = "lattice_riscv.v:50510.12-50510.59" *)
  wire [7:0] builder_csr_bankarray_interface3_bank_bus_dat_r_TMR_0;
  (* src = "lattice_riscv.v:50510.12-50510.59" *)
  wire [7:0] builder_csr_bankarray_interface3_bank_bus_dat_r_TMR_1;
  (* src = "lattice_riscv.v:50510.12-50510.59" *)
  wire [7:0] builder_csr_bankarray_interface3_bank_bus_dat_r_TMR_2;
  (* src = "lattice_riscv.v:51205.6-51205.36" *)
  wire builder_csr_bankarray_sel_r_QN;
  (* src = "lattice_riscv.v:50694.6-50694.33" *)
  wire builder_csr_bankarray_sel_r_TMR_0;
  (* src = "lattice_riscv.v:50694.6-50694.33" *)
  wire builder_csr_bankarray_sel_r_TMR_1;
  (* src = "lattice_riscv.v:50694.6-50694.33" *)
  wire builder_csr_bankarray_sel_r_TMR_2;
  (* src = "lattice_riscv.v:50728.6-50728.40" *)
  wire builder_csr_bankarray_sel_r_r_0_a2_TMR_0;
  (* src = "lattice_riscv.v:50728.6-50728.40" *)
  wire builder_csr_bankarray_sel_r_r_0_a2_TMR_1;
  (* src = "lattice_riscv.v:50728.6-50728.40" *)
  wire builder_csr_bankarray_sel_r_r_0_a2_TMR_2;
  (* src = "lattice_riscv.v:51206.6-51206.22" *)
  wire builder_grant_QN;
  (* src = "lattice_riscv.v:50671.6-50671.19" *)
  wire builder_grant_TMR_0;
  (* src = "lattice_riscv.v:50671.6-50671.19" *)
  wire builder_grant_TMR_1;
  (* src = "lattice_riscv.v:50671.6-50671.19" *)
  wire builder_grant_TMR_2;
  (* src = "lattice_riscv.v:51207.6-51207.27" *)
  wire builder_grant_fast_QN;
  (* src = "lattice_riscv.v:51177.6-51177.24" *)
  wire builder_grant_fast_TMR_0;
  (* src = "lattice_riscv.v:51177.6-51177.24" *)
  wire builder_grant_fast_TMR_1;
  (* src = "lattice_riscv.v:51177.6-51177.24" *)
  wire builder_grant_fast_TMR_2;
  (* src = "lattice_riscv.v:51208.6-51208.27" *)
  wire builder_grant_rep1_QN;
  (* src = "lattice_riscv.v:51179.6-51179.24" *)
  wire builder_grant_rep1_TMR_0;
  (* src = "lattice_riscv.v:51179.6-51179.24" *)
  wire builder_grant_rep1_TMR_1;
  (* src = "lattice_riscv.v:51179.6-51179.24" *)
  wire builder_grant_rep1_TMR_2;
  (* src = "lattice_riscv.v:51209.6-51209.27" *)
  wire builder_grant_rep2_QN;
  (* src = "lattice_riscv.v:51181.6-51181.24" *)
  wire builder_grant_rep2_TMR_0;
  (* src = "lattice_riscv.v:51181.6-51181.24" *)
  wire builder_grant_rep2_TMR_1;
  (* src = "lattice_riscv.v:51181.6-51181.24" *)
  wire builder_grant_rep2_TMR_2;
  (* src = "lattice_riscv.v:50677.6-50677.19" *)
  wire builder_regs0_TMR_0;
  (* src = "lattice_riscv.v:50677.6-50677.19" *)
  wire builder_regs0_TMR_1;
  (* src = "lattice_riscv.v:50677.6-50677.19" *)
  wire builder_regs0_TMR_2;
  (* src = "lattice_riscv.v:51210.6-51210.22" *)
  wire builder_regs1_QN;
  (* src = "lattice_riscv.v:50668.6-50668.19" *)
  wire builder_regs1_TMR_0;
  (* src = "lattice_riscv.v:50668.6-50668.19" *)
  wire builder_regs1_TMR_1;
  (* src = "lattice_riscv.v:50668.6-50668.19" *)
  wire builder_regs1_TMR_2;
  (* src = "lattice_riscv.v:50659.6-50659.19" *)
  wire builder_rst10_TMR_0;
  (* src = "lattice_riscv.v:50659.6-50659.19" *)
  wire builder_rst10_TMR_1;
  (* src = "lattice_riscv.v:50659.6-50659.19" *)
  wire builder_rst10_TMR_2;
  (* src = "lattice_riscv.v:50661.6-50661.19" *)
  wire builder_rst11_TMR_0;
  (* src = "lattice_riscv.v:50661.6-50661.19" *)
  wire builder_rst11_TMR_1;
  (* src = "lattice_riscv.v:50661.6-50661.19" *)
  wire builder_rst11_TMR_2;
  (* src = "lattice_riscv.v:50534.12-50534.31" *)
  wire builder_slave_sel_2_TMR_0;
  (* src = "lattice_riscv.v:50534.12-50534.31" *)
  wire builder_slave_sel_2_TMR_1;
  (* src = "lattice_riscv.v:50534.12-50534.31" *)
  wire builder_slave_sel_2_TMR_2;
  (* src = "lattice_riscv.v:50590.12-50590.34" *)
  wire [2:0] builder_slave_sel_r_QN;
  (* src = "lattice_riscv.v:50502.12-50502.31" *)
  wire [2:0] builder_slave_sel_r_TMR_0;
  (* src = "lattice_riscv.v:50502.12-50502.31" *)
  wire [2:0] builder_slave_sel_r_TMR_1;
  (* src = "lattice_riscv.v:50502.12-50502.31" *)
  wire [2:0] builder_slave_sel_r_TMR_2;
  (* src = "lattice_riscv.v:50528.12-50528.38" *)
  wire builder_slave_sel_r_r_0_a2_TMR_0;
  (* src = "lattice_riscv.v:50528.12-50528.38" *)
  wire builder_slave_sel_r_r_0_a2_TMR_1;
  (* src = "lattice_riscv.v:50528.12-50528.38" *)
  wire builder_slave_sel_r_r_0_a2_TMR_2;
  (* src = "lattice_riscv.v:50745.6-50745.18" *)
  wire builder_wait_TMR_0;
  (* src = "lattice_riscv.v:50745.6-50745.18" *)
  wire builder_wait_TMR_1;
  (* src = "lattice_riscv.v:50745.6-50745.18" *)
  wire builder_wait_TMR_2;
  (* src = "lattice_riscv.v:50508.13-50508.26" *)
  wire [30:0] dsp_join_kb_0_TMR_0;
  (* src = "lattice_riscv.v:50508.13-50508.26" *)
  wire [30:0] dsp_join_kb_0_TMR_1;
  (* src = "lattice_riscv.v:50508.13-50508.26" *)
  wire [30:0] dsp_join_kb_0_TMR_2;
  (* src = "lattice_riscv.v:50493.13-50493.27" *)
  wire [19:1] dsp_join_kb_25_TMR_0;
  (* src = "lattice_riscv.v:50493.13-50493.27" *)
  wire [19:1] dsp_join_kb_25_TMR_1;
  (* src = "lattice_riscv.v:50493.13-50493.27" *)
  wire [19:1] dsp_join_kb_25_TMR_2;
  (* src = "lattice_riscv.v:50625.14-50625.30" *)
  wire dsp_join_kb_25_i_TMR_0;
  (* src = "lattice_riscv.v:50625.14-50625.30" *)
  wire dsp_join_kb_25_i_TMR_1;
  (* src = "lattice_riscv.v:50625.14-50625.30" *)
  wire dsp_join_kb_25_i_TMR_2;
  (* src = "lattice_riscv.v:50516.13-50516.27" *)
  wire [31:0] dsp_join_kb_26_TMR_0;
  (* src = "lattice_riscv.v:50516.13-50516.27" *)
  wire [31:0] dsp_join_kb_26_TMR_1;
  (* src = "lattice_riscv.v:50516.13-50516.27" *)
  wire [31:0] dsp_join_kb_26_TMR_2;
  (* src = "lattice_riscv.v:50517.13-50517.27" *)
  wire [31:0] dsp_join_kb_27_TMR_0;
  (* src = "lattice_riscv.v:50517.13-50517.27" *)
  wire [31:0] dsp_join_kb_27_TMR_1;
  (* src = "lattice_riscv.v:50517.13-50517.27" *)
  wire [31:0] dsp_join_kb_27_TMR_2;
  (* src = "lattice_riscv.v:50536.13-50536.24" *)
  wire [30:0] dsp_join_kb_TMR_0;
  (* src = "lattice_riscv.v:50536.13-50536.24" *)
  wire [30:0] dsp_join_kb_TMR_1;
  (* src = "lattice_riscv.v:50536.13-50536.24" *)
  wire [30:0] dsp_join_kb_TMR_2;
  (* src = "lattice_riscv.v:50736.6-50736.20" *)
  wire dsp_split_kb_0_TMR_0;
  (* src = "lattice_riscv.v:50736.6-50736.20" *)
  wire dsp_split_kb_0_TMR_1;
  (* src = "lattice_riscv.v:50736.6-50736.20" *)
  wire dsp_split_kb_0_TMR_2;
  (* src = "lattice_riscv.v:50859.6-50859.20" *)
  wire dsp_split_kb_1_TMR_0;
  (* src = "lattice_riscv.v:50859.6-50859.20" *)
  wire dsp_split_kb_1_TMR_1;
  (* src = "lattice_riscv.v:50859.6-50859.20" *)
  wire dsp_split_kb_1_TMR_2;
  (* src = "lattice_riscv.v:50447.7-50447.11" *)
  input gsrn;
  wire gsrn;
  (* src = "lattice_riscv.v:51185.6-51185.12" *)
  wire gsrn_c;
  (* src = "lattice_riscv.v:51247.6-51247.14" *)
  wire gsrn_c_i_TMR_0;
  (* src = "lattice_riscv.v:51247.6-51247.14" *)
  wire gsrn_c_i_TMR_1;
  (* src = "lattice_riscv.v:51247.6-51247.14" *)
  wire gsrn_c_i_TMR_2;
  (* src = "lattice_riscv.v:51109.6-51109.9" *)
  wire m10_TMR_0;
  (* src = "lattice_riscv.v:51109.6-51109.9" *)
  wire m10_TMR_1;
  (* src = "lattice_riscv.v:51109.6-51109.9" *)
  wire m10_TMR_2;
  (* src = "lattice_riscv.v:51110.6-51110.9" *)
  wire m11_TMR_0;
  (* src = "lattice_riscv.v:51110.6-51110.9" *)
  wire m11_TMR_1;
  (* src = "lattice_riscv.v:51110.6-51110.9" *)
  wire m11_TMR_2;
  (* src = "lattice_riscv.v:51112.6-51112.9" *)
  wire m18_TMR_0;
  (* src = "lattice_riscv.v:51112.6-51112.9" *)
  wire m18_TMR_1;
  (* src = "lattice_riscv.v:51112.6-51112.9" *)
  wire m18_TMR_2;
  (* src = "lattice_riscv.v:51113.6-51113.9" *)
  wire m30_TMR_0;
  (* src = "lattice_riscv.v:51113.6-51113.9" *)
  wire m30_TMR_1;
  (* src = "lattice_riscv.v:51113.6-51113.9" *)
  wire m30_TMR_2;
  (* src = "lattice_riscv.v:51106.6-51106.8" *)
  wire m3_TMR_0;
  (* src = "lattice_riscv.v:51106.6-51106.8" *)
  wire m3_TMR_1;
  (* src = "lattice_riscv.v:51106.6-51106.8" *)
  wire m3_TMR_2;
  (* src = "lattice_riscv.v:51115.6-51115.9" *)
  wire m40_TMR_0;
  (* src = "lattice_riscv.v:51115.6-51115.9" *)
  wire m40_TMR_1;
  (* src = "lattice_riscv.v:51115.6-51115.9" *)
  wire m40_TMR_2;
  (* src = "lattice_riscv.v:51116.6-51116.9" *)
  wire m45_TMR_0;
  (* src = "lattice_riscv.v:51116.6-51116.9" *)
  wire m45_TMR_1;
  (* src = "lattice_riscv.v:51116.6-51116.9" *)
  wire m45_TMR_2;
  (* src = "lattice_riscv.v:51117.6-51117.9" *)
  wire m51_TMR_0;
  (* src = "lattice_riscv.v:51117.6-51117.9" *)
  wire m51_TMR_1;
  (* src = "lattice_riscv.v:51117.6-51117.9" *)
  wire m51_TMR_2;
  (* src = "lattice_riscv.v:51118.6-51118.9" *)
  wire m52_TMR_0;
  (* src = "lattice_riscv.v:51118.6-51118.9" *)
  wire m52_TMR_1;
  (* src = "lattice_riscv.v:51118.6-51118.9" *)
  wire m52_TMR_2;
  (* src = "lattice_riscv.v:51119.6-51119.9" *)
  wire m57_TMR_0;
  (* src = "lattice_riscv.v:51119.6-51119.9" *)
  wire m57_TMR_1;
  (* src = "lattice_riscv.v:51119.6-51119.9" *)
  wire m57_TMR_2;
  (* src = "lattice_riscv.v:51120.6-51120.9" *)
  wire m64_TMR_0;
  (* src = "lattice_riscv.v:51120.6-51120.9" *)
  wire m64_TMR_1;
  (* src = "lattice_riscv.v:51120.6-51120.9" *)
  wire m64_TMR_2;
  (* src = "lattice_riscv.v:51121.6-51121.9" *)
  wire m68_TMR_0;
  (* src = "lattice_riscv.v:51121.6-51121.9" *)
  wire m68_TMR_1;
  (* src = "lattice_riscv.v:51121.6-51121.9" *)
  wire m68_TMR_2;
  (* src = "lattice_riscv.v:51107.6-51107.8" *)
  wire m6_TMR_0;
  (* src = "lattice_riscv.v:51107.6-51107.8" *)
  wire m6_TMR_1;
  (* src = "lattice_riscv.v:51107.6-51107.8" *)
  wire m6_TMR_2;
  (* src = "lattice_riscv.v:51122.6-51122.9" *)
  wire m70_TMR_0;
  (* src = "lattice_riscv.v:51122.6-51122.9" *)
  wire m70_TMR_1;
  (* src = "lattice_riscv.v:51122.6-51122.9" *)
  wire m70_TMR_2;
  (* src = "lattice_riscv.v:51123.6-51123.9" *)
  wire m71_TMR_0;
  (* src = "lattice_riscv.v:51123.6-51123.9" *)
  wire m71_TMR_1;
  (* src = "lattice_riscv.v:51123.6-51123.9" *)
  wire m71_TMR_2;
  (* src = "lattice_riscv.v:51124.6-51124.9" *)
  wire m73_TMR_0;
  (* src = "lattice_riscv.v:51124.6-51124.9" *)
  wire m73_TMR_1;
  (* src = "lattice_riscv.v:51124.6-51124.9" *)
  wire m73_TMR_2;
  (* src = "lattice_riscv.v:51125.6-51125.9" *)
  wire m74_TMR_0;
  (* src = "lattice_riscv.v:51125.6-51125.9" *)
  wire m74_TMR_1;
  (* src = "lattice_riscv.v:51125.6-51125.9" *)
  wire m74_TMR_2;
  (* src = "lattice_riscv.v:51126.6-51126.9" *)
  wire m84_TMR_0;
  (* src = "lattice_riscv.v:51126.6-51126.9" *)
  wire m84_TMR_1;
  (* src = "lattice_riscv.v:51126.6-51126.9" *)
  wire m84_TMR_2;
  (* src = "lattice_riscv.v:51127.6-51127.9" *)
  wire m86_TMR_0;
  (* src = "lattice_riscv.v:51127.6-51127.9" *)
  wire m86_TMR_1;
  (* src = "lattice_riscv.v:51127.6-51127.9" *)
  wire m86_TMR_2;
  (* src = "lattice_riscv.v:51108.6-51108.8" *)
  wire m8_TMR_0;
  (* src = "lattice_riscv.v:51108.6-51108.8" *)
  wire m8_TMR_1;
  (* src = "lattice_riscv.v:51108.6-51108.8" *)
  wire m8_TMR_2;
  (* src = "lattice_riscv.v:50591.12-50591.44" *)
  wire main_basesoc_bus_errors_0_mod_QN;
  (* src = "lattice_riscv.v:50552.12-50552.45" *)
  wire main_basesoc_bus_errors_0_mod_RNO_TMR_0;
  (* src = "lattice_riscv.v:50552.12-50552.45" *)
  wire main_basesoc_bus_errors_0_mod_RNO_TMR_1;
  (* src = "lattice_riscv.v:50552.12-50552.45" *)
  wire main_basesoc_bus_errors_0_mod_RNO_TMR_2;
  (* src = "lattice_riscv.v:50698.6-50698.38" *)
  wire main_basesoc_bus_errors_0_sqmuxa_TMR_0;
  (* src = "lattice_riscv.v:50698.6-50698.38" *)
  wire main_basesoc_bus_errors_0_sqmuxa_TMR_1;
  (* src = "lattice_riscv.v:50698.6-50698.38" *)
  wire main_basesoc_bus_errors_0_sqmuxa_TMR_2;
  (* src = "lattice_riscv.v:50592.13-50592.43" *)
  wire [31:1] main_basesoc_bus_errors_mod_QN;
  (* src = "lattice_riscv.v:51211.6-51211.33" *)
  wire main_basesoc_ram_bus_ack_QN;
  (* src = "lattice_riscv.v:50672.6-50672.30" *)
  wire main_basesoc_ram_bus_ack_TMR_0;
  (* src = "lattice_riscv.v:50672.6-50672.30" *)
  wire main_basesoc_ram_bus_ack_TMR_1;
  (* src = "lattice_riscv.v:50672.6-50672.30" *)
  wire main_basesoc_ram_bus_ack_TMR_2;
  (* src = "lattice_riscv.v:50726.6-50726.32" *)
  wire main_basesoc_ram_bus_ack_r_TMR_0;
  (* src = "lattice_riscv.v:50726.6-50726.32" *)
  wire main_basesoc_ram_bus_ack_r_TMR_1;
  (* src = "lattice_riscv.v:50726.6-50726.32" *)
  wire main_basesoc_ram_bus_ack_r_TMR_2;
  (* src = "lattice_riscv.v:51212.6-51212.30" *)
  wire main_basesoc_reset_re_QN;
  (* src = "lattice_riscv.v:50691.6-50691.27" *)
  wire main_basesoc_reset_re_TMR_0;
  (* src = "lattice_riscv.v:50691.6-50691.27" *)
  wire main_basesoc_reset_re_TMR_1;
  (* src = "lattice_riscv.v:50691.6-50691.27" *)
  wire main_basesoc_reset_re_TMR_2;
  (* src = "lattice_riscv.v:50713.6-50713.41" *)
  wire main_basesoc_reset_storage_0_sqmuxa_TMR_0;
  (* src = "lattice_riscv.v:50713.6-50713.41" *)
  wire main_basesoc_reset_storage_0_sqmuxa_TMR_1;
  (* src = "lattice_riscv.v:50713.6-50713.41" *)
  wire main_basesoc_reset_storage_0_sqmuxa_TMR_2;
  (* src = "lattice_riscv.v:50593.12-50593.41" *)
  wire [1:0] main_basesoc_reset_storage_QN;
  (* src = "lattice_riscv.v:50503.12-50503.38" *)
  wire [1:0] main_basesoc_reset_storage_TMR_0;
  (* src = "lattice_riscv.v:50503.12-50503.38" *)
  wire [1:0] main_basesoc_reset_storage_TMR_1;
  (* src = "lattice_riscv.v:50503.12-50503.38" *)
  wire [1:0] main_basesoc_reset_storage_TMR_2;
  (* src = "lattice_riscv.v:51183.6-51183.34" *)
  wire \main_basesoc_rx_count_0_.fb_TMR_0 ;
  (* src = "lattice_riscv.v:51183.6-51183.34" *)
  wire \main_basesoc_rx_count_0_.fb_TMR_1 ;
  (* src = "lattice_riscv.v:51183.6-51183.34" *)
  wire \main_basesoc_rx_count_0_.fb_TMR_2 ;
  (* src = "lattice_riscv.v:50594.12-50594.36" *)
  wire [3:0] main_basesoc_rx_count_QN;
  (* src = "lattice_riscv.v:50491.12-50491.33" *)
  wire [3:1] main_basesoc_rx_count_TMR_0;
  (* src = "lattice_riscv.v:50491.12-50491.33" *)
  wire [3:1] main_basesoc_rx_count_TMR_1;
  (* src = "lattice_riscv.v:50491.12-50491.33" *)
  wire [3:1] main_basesoc_rx_count_TMR_2;
  (* src = "lattice_riscv.v:50533.12-50533.56" *)
  wire [3:1] main_basesoc_rx_count_rs232phyrx_next_value0_TMR_0;
  (* src = "lattice_riscv.v:50533.12-50533.56" *)
  wire [3:1] main_basesoc_rx_count_rs232phyrx_next_value0_TMR_1;
  (* src = "lattice_riscv.v:50533.12-50533.56" *)
  wire [3:1] main_basesoc_rx_count_rs232phyrx_next_value0_TMR_2;
  (* src = "lattice_riscv.v:50690.6-50690.53" *)
  wire main_basesoc_rx_count_rs232phyrx_next_value_ce0_TMR_0;
  (* src = "lattice_riscv.v:50690.6-50690.53" *)
  wire main_basesoc_rx_count_rs232phyrx_next_value_ce0_TMR_1;
  (* src = "lattice_riscv.v:50690.6-50690.53" *)
  wire main_basesoc_rx_count_rs232phyrx_next_value_ce0_TMR_2;
  (* src = "lattice_riscv.v:50595.12-50595.35" *)
  wire [7:0] main_basesoc_rx_data_QN;
  (* src = "lattice_riscv.v:50504.12-50504.32" *)
  wire [7:0] main_basesoc_rx_data_TMR_0;
  (* src = "lattice_riscv.v:50504.12-50504.32" *)
  wire [7:0] main_basesoc_rx_data_TMR_1;
  (* src = "lattice_riscv.v:50504.12-50504.32" *)
  wire [7:0] main_basesoc_rx_data_TMR_2;
  (* src = "lattice_riscv.v:50687.6-50687.58" *)
  wire main_basesoc_rx_data_rs232phyrx_next_value1_0_sqmuxa_TMR_0;
  (* src = "lattice_riscv.v:50687.6-50687.58" *)
  wire main_basesoc_rx_data_rs232phyrx_next_value1_0_sqmuxa_TMR_1;
  (* src = "lattice_riscv.v:50687.6-50687.58" *)
  wire main_basesoc_rx_data_rs232phyrx_next_value1_0_sqmuxa_TMR_2;
  (* src = "lattice_riscv.v:50596.14-50596.38" *)
  wire main_basesoc_rx_phase_QN;
  (* src = "lattice_riscv.v:50597.13-50597.41" *)
  wire [30:0] main_basesoc_rx_phase_mod_QN;
  (* src = "lattice_riscv.v:50550.12-50550.41" *)
  wire main_basesoc_rx_phase_mod_RNO_TMR_0;
  (* src = "lattice_riscv.v:50550.12-50550.41" *)
  wire main_basesoc_rx_phase_mod_RNO_TMR_1;
  (* src = "lattice_riscv.v:50550.12-50550.41" *)
  wire main_basesoc_rx_phase_mod_RNO_TMR_2;
  (* src = "lattice_riscv.v:51213.6-51213.29" *)
  wire main_basesoc_rx_rx_d_QN;
  (* src = "lattice_riscv.v:50689.6-50689.26" *)
  wire main_basesoc_rx_rx_d_TMR_0;
  (* src = "lattice_riscv.v:50689.6-50689.26" *)
  wire main_basesoc_rx_rx_d_TMR_1;
  (* src = "lattice_riscv.v:50689.6-50689.26" *)
  wire main_basesoc_rx_rx_d_TMR_2;
  (* src = "lattice_riscv.v:50511.12-50511.47" *)
  wire [7:0] main_basesoc_rx_source_payload_data_TMR_0;
  (* src = "lattice_riscv.v:50511.12-50511.47" *)
  wire [7:0] main_basesoc_rx_source_payload_data_TMR_1;
  (* src = "lattice_riscv.v:50511.12-50511.47" *)
  wire [7:0] main_basesoc_rx_source_payload_data_TMR_2;
  (* src = "lattice_riscv.v:50730.6-50730.28" *)
  wire main_basesoc_rx_tick_0_TMR_0;
  (* src = "lattice_riscv.v:50730.6-50730.28" *)
  wire main_basesoc_rx_tick_0_TMR_1;
  (* src = "lattice_riscv.v:50730.6-50730.28" *)
  wire main_basesoc_rx_tick_0_TMR_2;
  (* src = "lattice_riscv.v:51214.6-51214.29" *)
  wire main_basesoc_rx_tick_QN;
  (* src = "lattice_riscv.v:50688.6-50688.26" *)
  wire main_basesoc_rx_tick_TMR_0;
  (* src = "lattice_riscv.v:50688.6-50688.26" *)
  wire main_basesoc_rx_tick_TMR_1;
  (* src = "lattice_riscv.v:50688.6-50688.26" *)
  wire main_basesoc_rx_tick_TMR_2;
  (* src = "lattice_riscv.v:50598.13-50598.44" *)
  wire [31:0] main_basesoc_scratch_storage_QN;
  (* src = "lattice_riscv.v:50522.13-50522.41" *)
  wire [31:0] main_basesoc_scratch_storage_TMR_0;
  (* src = "lattice_riscv.v:50522.13-50522.41" *)
  wire [31:0] main_basesoc_scratch_storage_TMR_1;
  (* src = "lattice_riscv.v:50522.13-50522.41" *)
  wire [31:0] main_basesoc_scratch_storage_TMR_2;
  (* src = "lattice_riscv.v:51103.6-51103.62" *)
  wire main_basesoc_serial_tx_rs232phytx_next_value1_1_sqmuxa_i_TMR_0;
  (* src = "lattice_riscv.v:51103.6-51103.62" *)
  wire main_basesoc_serial_tx_rs232phytx_next_value1_1_sqmuxa_i_TMR_1;
  (* src = "lattice_riscv.v:51103.6-51103.62" *)
  wire main_basesoc_serial_tx_rs232phytx_next_value1_1_sqmuxa_i_TMR_2;
  (* src = "lattice_riscv.v:51215.6-51215.38" *)
  wire main_basesoc_timer_en_storage_QN;
  (* src = "lattice_riscv.v:50665.6-50665.35" *)
  wire main_basesoc_timer_en_storage_TMR_0;
  (* src = "lattice_riscv.v:50665.6-50665.35" *)
  wire main_basesoc_timer_en_storage_TMR_1;
  (* src = "lattice_riscv.v:50665.6-50665.35" *)
  wire main_basesoc_timer_en_storage_TMR_2;
  (* src = "lattice_riscv.v:51216.6-51216.42" *)
  wire main_basesoc_timer_enable_storage_QN;
  (* src = "lattice_riscv.v:50685.6-50685.39" *)
  wire main_basesoc_timer_enable_storage_TMR_0;
  (* src = "lattice_riscv.v:50685.6-50685.39" *)
  wire main_basesoc_timer_enable_storage_TMR_1;
  (* src = "lattice_riscv.v:50685.6-50685.39" *)
  wire main_basesoc_timer_enable_storage_TMR_2;
  (* src = "lattice_riscv.v:50599.13-50599.53" *)
  wire [30:0] main_basesoc_timer_load_storage_0_mod_QN;
  (* src = "lattice_riscv.v:50551.12-50551.53" *)
  wire main_basesoc_timer_load_storage_0_mod_RNO_TMR_0;
  (* src = "lattice_riscv.v:50551.12-50551.53" *)
  wire main_basesoc_timer_load_storage_0_mod_RNO_TMR_1;
  (* src = "lattice_riscv.v:50551.12-50551.53" *)
  wire main_basesoc_timer_load_storage_0_mod_RNO_TMR_2;
  (* src = "lattice_riscv.v:50600.13-50600.51" *)
  wire [31:1] main_basesoc_timer_load_storage_mod_QN;
  (* src = "lattice_riscv.v:50716.6-50716.43" *)
  wire main_basesoc_timer_pending_r_0_sqmuxa_TMR_0;
  (* src = "lattice_riscv.v:50716.6-50716.43" *)
  wire main_basesoc_timer_pending_r_0_sqmuxa_TMR_1;
  (* src = "lattice_riscv.v:50716.6-50716.43" *)
  wire main_basesoc_timer_pending_r_0_sqmuxa_TMR_2;
  (* src = "lattice_riscv.v:51217.6-51217.37" *)
  wire main_basesoc_timer_pending_r_QN;
  (* src = "lattice_riscv.v:50683.6-50683.34" *)
  wire main_basesoc_timer_pending_r_TMR_0;
  (* src = "lattice_riscv.v:50683.6-50683.34" *)
  wire main_basesoc_timer_pending_r_TMR_1;
  (* src = "lattice_riscv.v:50683.6-50683.34" *)
  wire main_basesoc_timer_pending_r_TMR_2;
  (* src = "lattice_riscv.v:51218.6-51218.38" *)
  wire main_basesoc_timer_pending_re_QN;
  (* src = "lattice_riscv.v:50682.6-50682.35" *)
  wire main_basesoc_timer_pending_re_TMR_0;
  (* src = "lattice_riscv.v:50682.6-50682.35" *)
  wire main_basesoc_timer_pending_re_TMR_1;
  (* src = "lattice_riscv.v:50682.6-50682.35" *)
  wire main_basesoc_timer_pending_re_TMR_2;
  (* src = "lattice_riscv.v:50601.13-50601.49" *)
  wire [31:0] main_basesoc_timer_reload_storage_QN;
  (* src = "lattice_riscv.v:50519.13-50519.46" *)
  wire [31:0] main_basesoc_timer_reload_storage_TMR_0;
  (* src = "lattice_riscv.v:50519.13-50519.46" *)
  wire [31:0] main_basesoc_timer_reload_storage_TMR_1;
  (* src = "lattice_riscv.v:50519.13-50519.46" *)
  wire [31:0] main_basesoc_timer_reload_storage_TMR_2;
  (* src = "lattice_riscv.v:51219.6-51219.43" *)
  wire main_basesoc_timer_update_value_re_QN;
  (* src = "lattice_riscv.v:50719.6-50719.40" *)
  wire main_basesoc_timer_update_value_re_TMR_0;
  (* src = "lattice_riscv.v:50719.6-50719.40" *)
  wire main_basesoc_timer_update_value_re_TMR_1;
  (* src = "lattice_riscv.v:50719.6-50719.40" *)
  wire main_basesoc_timer_update_value_re_TMR_2;
  (* src = "lattice_riscv.v:50715.6-50715.54" *)
  wire main_basesoc_timer_update_value_storage_0_sqmuxa_TMR_0;
  (* src = "lattice_riscv.v:50715.6-50715.54" *)
  wire main_basesoc_timer_update_value_storage_0_sqmuxa_TMR_1;
  (* src = "lattice_riscv.v:50715.6-50715.54" *)
  wire main_basesoc_timer_update_value_storage_0_sqmuxa_TMR_2;
  (* src = "lattice_riscv.v:51220.6-51220.48" *)
  wire main_basesoc_timer_update_value_storage_QN;
  (* src = "lattice_riscv.v:50712.6-50712.45" *)
  wire main_basesoc_timer_update_value_storage_TMR_0;
  (* src = "lattice_riscv.v:50712.6-50712.45" *)
  wire main_basesoc_timer_update_value_storage_TMR_1;
  (* src = "lattice_riscv.v:50712.6-50712.45" *)
  wire main_basesoc_timer_update_value_storage_TMR_2;
  (* src = "lattice_riscv.v:50602.13-50602.46" *)
  wire [31:0] main_basesoc_timer_value_0_mod_QN;
  (* src = "lattice_riscv.v:50546.12-50546.46" *)
  wire main_basesoc_timer_value_0_mod_RNO_TMR_0;
  (* src = "lattice_riscv.v:50546.12-50546.46" *)
  wire main_basesoc_timer_value_0_mod_RNO_TMR_1;
  (* src = "lattice_riscv.v:50546.12-50546.46" *)
  wire main_basesoc_timer_value_0_mod_RNO_TMR_2;
  (* src = "lattice_riscv.v:50603.13-50603.47" *)
  wire [31:0] main_basesoc_timer_value_status_QN;
  (* src = "lattice_riscv.v:50525.13-50525.44" *)
  wire [31:0] main_basesoc_timer_value_status_TMR_0;
  (* src = "lattice_riscv.v:50525.13-50525.44" *)
  wire [31:0] main_basesoc_timer_value_status_TMR_1;
  (* src = "lattice_riscv.v:50525.13-50525.44" *)
  wire [31:0] main_basesoc_timer_value_status_TMR_2;
  (* src = "lattice_riscv.v:51221.6-51221.40" *)
  wire main_basesoc_timer_zero_pending_QN;
  (* src = "lattice_riscv.v:50684.6-50684.37" *)
  wire main_basesoc_timer_zero_pending_TMR_0;
  (* src = "lattice_riscv.v:50684.6-50684.37" *)
  wire main_basesoc_timer_zero_pending_TMR_1;
  (* src = "lattice_riscv.v:50684.6-50684.37" *)
  wire main_basesoc_timer_zero_pending_TMR_2;
  (* src = "lattice_riscv.v:50735.6-50735.37" *)
  wire main_basesoc_timer_zero_trigger_TMR_0;
  (* src = "lattice_riscv.v:50735.6-50735.37" *)
  wire main_basesoc_timer_zero_trigger_TMR_1;
  (* src = "lattice_riscv.v:50735.6-50735.37" *)
  wire main_basesoc_timer_zero_trigger_TMR_2;
  (* src = "lattice_riscv.v:51222.6-51222.42" *)
  wire main_basesoc_timer_zero_trigger_d_QN;
  (* src = "lattice_riscv.v:50675.6-50675.39" *)
  wire main_basesoc_timer_zero_trigger_d_TMR_0;
  (* src = "lattice_riscv.v:50675.6-50675.39" *)
  wire main_basesoc_timer_zero_trigger_d_TMR_1;
  (* src = "lattice_riscv.v:50675.6-50675.39" *)
  wire main_basesoc_timer_zero_trigger_d_TMR_2;
  (* src = "lattice_riscv.v:51184.6-51184.34" *)
  wire \main_basesoc_tx_count_0_.fb_TMR_0 ;
  (* src = "lattice_riscv.v:51184.6-51184.34" *)
  wire \main_basesoc_tx_count_0_.fb_TMR_1 ;
  (* src = "lattice_riscv.v:51184.6-51184.34" *)
  wire \main_basesoc_tx_count_0_.fb_TMR_2 ;
  (* src = "lattice_riscv.v:50604.12-50604.36" *)
  wire [3:0] main_basesoc_tx_count_QN;
  (* src = "lattice_riscv.v:50490.12-50490.33" *)
  wire [3:1] main_basesoc_tx_count_TMR_0;
  (* src = "lattice_riscv.v:50490.12-50490.33" *)
  wire [3:1] main_basesoc_tx_count_TMR_1;
  (* src = "lattice_riscv.v:50490.12-50490.33" *)
  wire [3:1] main_basesoc_tx_count_TMR_2;
  (* src = "lattice_riscv.v:50535.12-50535.56" *)
  wire [3:1] main_basesoc_tx_count_rs232phytx_next_value0_TMR_0;
  (* src = "lattice_riscv.v:50535.12-50535.56" *)
  wire [3:1] main_basesoc_tx_count_rs232phytx_next_value0_TMR_1;
  (* src = "lattice_riscv.v:50535.12-50535.56" *)
  wire [3:1] main_basesoc_tx_count_rs232phytx_next_value0_TMR_2;
  (* src = "lattice_riscv.v:50605.12-50605.35" *)
  wire [7:0] main_basesoc_tx_data_QN;
  (* src = "lattice_riscv.v:50507.12-50507.32" *)
  wire [7:0] main_basesoc_tx_data_TMR_0;
  (* src = "lattice_riscv.v:50507.12-50507.32" *)
  wire [7:0] main_basesoc_tx_data_TMR_1;
  (* src = "lattice_riscv.v:50507.12-50507.32" *)
  wire [7:0] main_basesoc_tx_data_TMR_2;
  (* src = "lattice_riscv.v:50746.6-50746.58" *)
  wire main_basesoc_tx_data_rs232phytx_next_value2_0_sqmuxa_TMR_0;
  (* src = "lattice_riscv.v:50746.6-50746.58" *)
  wire main_basesoc_tx_data_rs232phytx_next_value2_0_sqmuxa_TMR_1;
  (* src = "lattice_riscv.v:50746.6-50746.58" *)
  wire main_basesoc_tx_data_rs232phytx_next_value2_0_sqmuxa_TMR_2;
  (* src = "lattice_riscv.v:50505.12-50505.55" *)
  wire [7:0] main_basesoc_tx_data_rs232phytx_next_value2_TMR_0;
  (* src = "lattice_riscv.v:50505.12-50505.55" *)
  wire [7:0] main_basesoc_tx_data_rs232phytx_next_value2_TMR_1;
  (* src = "lattice_riscv.v:50505.12-50505.55" *)
  wire [7:0] main_basesoc_tx_data_rs232phytx_next_value2_TMR_2;
  (* src = "lattice_riscv.v:50678.6-50678.54" *)
  wire main_basesoc_tx_data_rs232phytx_next_value_ce2_1_TMR_0;
  (* src = "lattice_riscv.v:50678.6-50678.54" *)
  wire main_basesoc_tx_data_rs232phytx_next_value_ce2_1_TMR_1;
  (* src = "lattice_riscv.v:50678.6-50678.54" *)
  wire main_basesoc_tx_data_rs232phytx_next_value_ce2_1_TMR_2;
  (* src = "lattice_riscv.v:50606.13-50606.37" *)
  wire [31:1] main_basesoc_tx_phase_QN;
  (* src = "lattice_riscv.v:50607.12-50607.40" *)
  wire main_basesoc_tx_phase_mod_QN;
  (* src = "lattice_riscv.v:50549.12-50549.41" *)
  wire main_basesoc_tx_phase_mod_RNO_TMR_0;
  (* src = "lattice_riscv.v:50549.12-50549.41" *)
  wire main_basesoc_tx_phase_mod_RNO_TMR_1;
  (* src = "lattice_riscv.v:50549.12-50549.41" *)
  wire main_basesoc_tx_phase_mod_RNO_TMR_2;
  (* src = "lattice_riscv.v:50729.6-50729.28" *)
  wire main_basesoc_tx_tick_0_TMR_0;
  (* src = "lattice_riscv.v:50729.6-50729.28" *)
  wire main_basesoc_tx_tick_0_TMR_1;
  (* src = "lattice_riscv.v:50729.6-50729.28" *)
  wire main_basesoc_tx_tick_0_TMR_2;
  (* src = "lattice_riscv.v:51223.6-51223.29" *)
  wire main_basesoc_tx_tick_QN;
  (* src = "lattice_riscv.v:50664.6-50664.26" *)
  wire main_basesoc_tx_tick_TMR_0;
  (* src = "lattice_riscv.v:50664.6-50664.26" *)
  wire main_basesoc_tx_tick_TMR_1;
  (* src = "lattice_riscv.v:50664.6-50664.26" *)
  wire main_basesoc_tx_tick_TMR_2;
  (* src = "lattice_riscv.v:50608.12-50608.47" *)
  wire [1:0] main_basesoc_uart_enable_storage_QN;
  (* src = "lattice_riscv.v:50497.12-50497.44" *)
  wire [1:0] main_basesoc_uart_enable_storage_TMR_0;
  (* src = "lattice_riscv.v:50497.12-50497.44" *)
  wire [1:0] main_basesoc_uart_enable_storage_TMR_1;
  (* src = "lattice_riscv.v:50497.12-50497.44" *)
  wire [1:0] main_basesoc_uart_enable_storage_TMR_2;
  (* src = "lattice_riscv.v:50717.6-50717.42" *)
  wire main_basesoc_uart_pending_r_0_sqmuxa_TMR_0;
  (* src = "lattice_riscv.v:50717.6-50717.42" *)
  wire main_basesoc_uart_pending_r_0_sqmuxa_TMR_1;
  (* src = "lattice_riscv.v:50717.6-50717.42" *)
  wire main_basesoc_uart_pending_r_0_sqmuxa_TMR_2;
  (* src = "lattice_riscv.v:50609.12-50609.42" *)
  wire [1:0] main_basesoc_uart_pending_r_QN;
  (* src = "lattice_riscv.v:50496.12-50496.39" *)
  wire [1:0] main_basesoc_uart_pending_r_TMR_0;
  (* src = "lattice_riscv.v:50496.12-50496.39" *)
  wire [1:0] main_basesoc_uart_pending_r_TMR_1;
  (* src = "lattice_riscv.v:50496.12-50496.39" *)
  wire [1:0] main_basesoc_uart_pending_r_TMR_2;
  (* src = "lattice_riscv.v:51224.6-51224.37" *)
  wire main_basesoc_uart_pending_re_QN;
  (* src = "lattice_riscv.v:50679.6-50679.34" *)
  wire main_basesoc_uart_pending_re_TMR_0;
  (* src = "lattice_riscv.v:50679.6-50679.34" *)
  wire main_basesoc_uart_pending_re_TMR_1;
  (* src = "lattice_riscv.v:50679.6-50679.34" *)
  wire main_basesoc_uart_pending_re_TMR_2;
  (* src = "lattice_riscv.v:50610.12-50610.48" *)
  wire [3:0] main_basesoc_uart_rx_fifo_consume_QN;
  (* src = "lattice_riscv.v:50559.12-50559.49" *)
  wire main_basesoc_uart_rx_fifo_consume_RNO_TMR_0;
  (* src = "lattice_riscv.v:50559.12-50559.49" *)
  wire main_basesoc_uart_rx_fifo_consume_RNO_TMR_1;
  (* src = "lattice_riscv.v:50559.12-50559.49" *)
  wire main_basesoc_uart_rx_fifo_consume_RNO_TMR_2;
  (* src = "lattice_riscv.v:50513.12-50513.45" *)
  wire [3:0] main_basesoc_uart_rx_fifo_consume_TMR_0;
  (* src = "lattice_riscv.v:50513.12-50513.45" *)
  wire [3:0] main_basesoc_uart_rx_fifo_consume_TMR_1;
  (* src = "lattice_riscv.v:50513.12-50513.45" *)
  wire [3:0] main_basesoc_uart_rx_fifo_consume_TMR_2;
  (* src = "lattice_riscv.v:50611.12-50611.53" *)
  wire [4:0] main_basesoc_uart_rx_fifo_level0_0_mod_QN;
  (* src = "lattice_riscv.v:50553.12-50553.54" *)
  wire main_basesoc_uart_rx_fifo_level0_0_mod_RNO_TMR_0;
  (* src = "lattice_riscv.v:50553.12-50553.54" *)
  wire main_basesoc_uart_rx_fifo_level0_0_mod_RNO_TMR_1;
  (* src = "lattice_riscv.v:50553.12-50553.54" *)
  wire main_basesoc_uart_rx_fifo_level0_0_mod_RNO_TMR_2;
  (* src = "lattice_riscv.v:50612.12-50612.51" *)
  wire [3:1] main_basesoc_uart_rx_fifo_level0_mod_QN;
  (* src = "lattice_riscv.v:50613.12-50613.48" *)
  wire [3:0] main_basesoc_uart_rx_fifo_produce_QN;
  (* src = "lattice_riscv.v:50561.12-50561.49" *)
  wire main_basesoc_uart_rx_fifo_produce_RNO_TMR_0;
  (* src = "lattice_riscv.v:50561.12-50561.49" *)
  wire main_basesoc_uart_rx_fifo_produce_RNO_TMR_1;
  (* src = "lattice_riscv.v:50561.12-50561.49" *)
  wire main_basesoc_uart_rx_fifo_produce_RNO_TMR_2;
  (* src = "lattice_riscv.v:50514.12-50514.45" *)
  wire [3:0] main_basesoc_uart_rx_fifo_produce_TMR_0;
  (* src = "lattice_riscv.v:50514.12-50514.45" *)
  wire [3:0] main_basesoc_uart_rx_fifo_produce_TMR_1;
  (* src = "lattice_riscv.v:50514.12-50514.45" *)
  wire [3:0] main_basesoc_uart_rx_fifo_produce_TMR_2;
  (* src = "lattice_riscv.v:51225.6-51225.43" *)
  wire main_basesoc_uart_rx_fifo_readable_QN;
  (* src = "lattice_riscv.v:50669.6-50669.40" *)
  wire main_basesoc_uart_rx_fifo_readable_TMR_0;
  (* src = "lattice_riscv.v:50669.6-50669.40" *)
  wire main_basesoc_uart_rx_fifo_readable_TMR_1;
  (* src = "lattice_riscv.v:50669.6-50669.40" *)
  wire main_basesoc_uart_rx_fifo_readable_TMR_2;
  (* src = "lattice_riscv.v:50696.6-50696.43" *)
  wire main_basesoc_uart_rx_fifo_syncfifo_re_TMR_0;
  (* src = "lattice_riscv.v:50696.6-50696.43" *)
  wire main_basesoc_uart_rx_fifo_syncfifo_re_TMR_1;
  (* src = "lattice_riscv.v:50696.6-50696.43" *)
  wire main_basesoc_uart_rx_fifo_syncfifo_re_TMR_2;
  (* src = "lattice_riscv.v:50700.6-50700.41" *)
  wire main_basesoc_uart_rx_fifo_wrport_we_TMR_0;
  (* src = "lattice_riscv.v:50700.6-50700.41" *)
  wire main_basesoc_uart_rx_fifo_wrport_we_TMR_1;
  (* src = "lattice_riscv.v:50700.6-50700.41" *)
  wire main_basesoc_uart_rx_fifo_wrport_we_TMR_2;
  (* src = "lattice_riscv.v:51226.6-51226.37" *)
  wire main_basesoc_uart_rx_pending_QN;
  (* src = "lattice_riscv.v:50681.6-50681.34" *)
  wire main_basesoc_uart_rx_pending_TMR_0;
  (* src = "lattice_riscv.v:50681.6-50681.34" *)
  wire main_basesoc_uart_rx_pending_TMR_1;
  (* src = "lattice_riscv.v:50681.6-50681.34" *)
  wire main_basesoc_uart_rx_pending_TMR_2;
  (* src = "lattice_riscv.v:51227.6-51227.39" *)
  wire main_basesoc_uart_rx_trigger_d_QN;
  (* src = "lattice_riscv.v:50674.6-50674.36" *)
  wire main_basesoc_uart_rx_trigger_d_TMR_0;
  (* src = "lattice_riscv.v:50674.6-50674.36" *)
  wire main_basesoc_uart_rx_trigger_d_TMR_1;
  (* src = "lattice_riscv.v:50674.6-50674.36" *)
  wire main_basesoc_uart_rx_trigger_d_TMR_2;
  (* src = "lattice_riscv.v:50614.12-50614.48" *)
  wire [3:0] main_basesoc_uart_tx_fifo_consume_QN;
  (* src = "lattice_riscv.v:50560.12-50560.49" *)
  wire main_basesoc_uart_tx_fifo_consume_RNO_TMR_0;
  (* src = "lattice_riscv.v:50560.12-50560.49" *)
  wire main_basesoc_uart_tx_fifo_consume_RNO_TMR_1;
  (* src = "lattice_riscv.v:50560.12-50560.49" *)
  wire main_basesoc_uart_tx_fifo_consume_RNO_TMR_2;
  (* src = "lattice_riscv.v:50518.12-50518.45" *)
  wire [3:0] main_basesoc_uart_tx_fifo_consume_TMR_0;
  (* src = "lattice_riscv.v:50518.12-50518.45" *)
  wire [3:0] main_basesoc_uart_tx_fifo_consume_TMR_1;
  (* src = "lattice_riscv.v:50518.12-50518.45" *)
  wire [3:0] main_basesoc_uart_tx_fifo_consume_TMR_2;
  (* src = "lattice_riscv.v:50615.12-50615.53" *)
  wire [4:0] main_basesoc_uart_tx_fifo_level0_0_mod_QN;
  (* src = "lattice_riscv.v:50582.12-50582.58" *)
  wire main_basesoc_uart_tx_fifo_level0_0_mod_RNIG0F3_TMR_0;
  (* src = "lattice_riscv.v:50582.12-50582.58" *)
  wire main_basesoc_uart_tx_fifo_level0_0_mod_RNIG0F3_TMR_1;
  (* src = "lattice_riscv.v:50582.12-50582.58" *)
  wire main_basesoc_uart_tx_fifo_level0_0_mod_RNIG0F3_TMR_2;
  (* src = "lattice_riscv.v:50554.12-50554.54" *)
  wire main_basesoc_uart_tx_fifo_level0_0_mod_RNO_TMR_0;
  (* src = "lattice_riscv.v:50554.12-50554.54" *)
  wire main_basesoc_uart_tx_fifo_level0_0_mod_RNO_TMR_1;
  (* src = "lattice_riscv.v:50554.12-50554.54" *)
  wire main_basesoc_uart_tx_fifo_level0_0_mod_RNO_TMR_2;
  (* src = "lattice_riscv.v:50616.12-50616.51" *)
  wire [3:1] main_basesoc_uart_tx_fifo_level0_mod_QN;
  (* src = "lattice_riscv.v:50617.12-50617.48" *)
  wire [3:0] main_basesoc_uart_tx_fifo_produce_QN;
  (* src = "lattice_riscv.v:50562.12-50562.49" *)
  wire main_basesoc_uart_tx_fifo_produce_RNO_TMR_0;
  (* src = "lattice_riscv.v:50562.12-50562.49" *)
  wire main_basesoc_uart_tx_fifo_produce_RNO_TMR_1;
  (* src = "lattice_riscv.v:50562.12-50562.49" *)
  wire main_basesoc_uart_tx_fifo_produce_RNO_TMR_2;
  (* src = "lattice_riscv.v:50524.12-50524.45" *)
  wire [3:0] main_basesoc_uart_tx_fifo_produce_TMR_0;
  (* src = "lattice_riscv.v:50524.12-50524.45" *)
  wire [3:0] main_basesoc_uart_tx_fifo_produce_TMR_1;
  (* src = "lattice_riscv.v:50524.12-50524.45" *)
  wire [3:0] main_basesoc_uart_tx_fifo_produce_TMR_2;
  (* src = "lattice_riscv.v:51228.6-51228.43" *)
  wire main_basesoc_uart_tx_fifo_readable_QN;
  (* src = "lattice_riscv.v:50663.6-50663.40" *)
  wire main_basesoc_uart_tx_fifo_readable_TMR_0;
  (* src = "lattice_riscv.v:50663.6-50663.40" *)
  wire main_basesoc_uart_tx_fifo_readable_TMR_1;
  (* src = "lattice_riscv.v:50663.6-50663.40" *)
  wire main_basesoc_uart_tx_fifo_readable_TMR_2;
  (* src = "lattice_riscv.v:50699.6-50699.43" *)
  wire main_basesoc_uart_tx_fifo_syncfifo_re_TMR_0;
  (* src = "lattice_riscv.v:50699.6-50699.43" *)
  wire main_basesoc_uart_tx_fifo_syncfifo_re_TMR_1;
  (* src = "lattice_riscv.v:50699.6-50699.43" *)
  wire main_basesoc_uart_tx_fifo_syncfifo_re_TMR_2;
  (* src = "lattice_riscv.v:50718.6-50718.41" *)
  wire main_basesoc_uart_tx_fifo_wrport_we_TMR_0;
  (* src = "lattice_riscv.v:50718.6-50718.41" *)
  wire main_basesoc_uart_tx_fifo_wrport_we_TMR_1;
  (* src = "lattice_riscv.v:50718.6-50718.41" *)
  wire main_basesoc_uart_tx_fifo_wrport_we_TMR_2;
  (* src = "lattice_riscv.v:51229.6-51229.37" *)
  wire main_basesoc_uart_tx_pending_QN;
  (* src = "lattice_riscv.v:50680.6-50680.34" *)
  wire main_basesoc_uart_tx_pending_TMR_0;
  (* src = "lattice_riscv.v:50680.6-50680.34" *)
  wire main_basesoc_uart_tx_pending_TMR_1;
  (* src = "lattice_riscv.v:50680.6-50680.34" *)
  wire main_basesoc_uart_tx_pending_TMR_2;
  (* src = "lattice_riscv.v:51230.6-51230.39" *)
  wire main_basesoc_uart_tx_trigger_d_QN;
  (* src = "lattice_riscv.v:50673.6-50673.36" *)
  wire main_basesoc_uart_tx_trigger_d_TMR_0;
  (* src = "lattice_riscv.v:50673.6-50673.36" *)
  wire main_basesoc_uart_tx_trigger_d_TMR_1;
  (* src = "lattice_riscv.v:50673.6-50673.36" *)
  wire main_basesoc_uart_tx_trigger_d_TMR_2;
  (* src = "lattice_riscv.v:51231.6-51231.21" *)
  wire main_bus_ack_QN;
  (* src = "lattice_riscv.v:50676.6-50676.18" *)
  wire main_bus_ack_TMR_0;
  (* src = "lattice_riscv.v:50676.6-50676.18" *)
  wire main_bus_ack_TMR_1;
  (* src = "lattice_riscv.v:50676.6-50676.18" *)
  wire main_bus_ack_TMR_2;
  (* src = "lattice_riscv.v:50727.6-50727.25" *)
  wire main_bus_ack_r_0_a2_TMR_0;
  (* src = "lattice_riscv.v:50727.6-50727.25" *)
  wire main_bus_ack_r_0_a2_TMR_1;
  (* src = "lattice_riscv.v:50727.6-50727.25" *)
  wire main_bus_ack_r_0_a2_TMR_2;
  (* src = "lattice_riscv.v:50618.13-50618.27" *)
  wire [13:0] main_chaser_QN;
  (* src = "lattice_riscv.v:50494.13-50494.24" *)
  wire [13:0] main_chaser_TMR_0;
  (* src = "lattice_riscv.v:50494.13-50494.24" *)
  wire [13:0] main_chaser_TMR_1;
  (* src = "lattice_riscv.v:50494.13-50494.24" *)
  wire [13:0] main_chaser_TMR_2;
  (* src = "lattice_riscv.v:50626.14-50626.27" *)
  wire main_chaser_i_TMR_0;
  (* src = "lattice_riscv.v:50626.14-50626.27" *)
  wire main_chaser_i_TMR_1;
  (* src = "lattice_riscv.v:50626.14-50626.27" *)
  wire main_chaser_i_TMR_2;
  (* src = "lattice_riscv.v:50986.6-50986.18" *)
  wire main_count_1_TMR_0;
  (* src = "lattice_riscv.v:50986.6-50986.18" *)
  wire main_count_1_TMR_1;
  (* src = "lattice_riscv.v:50986.6-50986.18" *)
  wire main_count_1_TMR_2;
  (* src = "lattice_riscv.v:51154.6-51154.29" *)
  wire main_count_1_cry_0_0_S0_TMR_0;
  (* src = "lattice_riscv.v:51154.6-51154.29" *)
  wire main_count_1_cry_0_0_S0_TMR_1;
  (* src = "lattice_riscv.v:51154.6-51154.29" *)
  wire main_count_1_cry_0_0_S0_TMR_2;
  (* src = "lattice_riscv.v:51148.6-51148.29" *)
  wire main_count_1_cry_0_0_S1_TMR_0;
  (* src = "lattice_riscv.v:51148.6-51148.29" *)
  wire main_count_1_cry_0_0_S1_TMR_1;
  (* src = "lattice_riscv.v:51148.6-51148.29" *)
  wire main_count_1_cry_0_0_S1_TMR_2;
  (* src = "lattice_riscv.v:51061.6-51061.24" *)
  wire main_count_1_cry_0_TMR_0;
  (* src = "lattice_riscv.v:51061.6-51061.24" *)
  wire main_count_1_cry_0_TMR_1;
  (* src = "lattice_riscv.v:51061.6-51061.24" *)
  wire main_count_1_cry_0_TMR_2;
  (* src = "lattice_riscv.v:51066.6-51066.25" *)
  wire main_count_1_cry_10_TMR_0;
  (* src = "lattice_riscv.v:51066.6-51066.25" *)
  wire main_count_1_cry_10_TMR_1;
  (* src = "lattice_riscv.v:51066.6-51066.25" *)
  wire main_count_1_cry_10_TMR_2;
  (* src = "lattice_riscv.v:50757.6-50757.30" *)
  wire main_count_1_cry_11_0_S0_TMR_0;
  (* src = "lattice_riscv.v:50757.6-50757.30" *)
  wire main_count_1_cry_11_0_S0_TMR_1;
  (* src = "lattice_riscv.v:50757.6-50757.30" *)
  wire main_count_1_cry_11_0_S0_TMR_2;
  (* src = "lattice_riscv.v:50758.6-50758.30" *)
  wire main_count_1_cry_11_0_S1_TMR_0;
  (* src = "lattice_riscv.v:50758.6-50758.30" *)
  wire main_count_1_cry_11_0_S1_TMR_1;
  (* src = "lattice_riscv.v:50758.6-50758.30" *)
  wire main_count_1_cry_11_0_S1_TMR_2;
  (* src = "lattice_riscv.v:51067.6-51067.25" *)
  wire main_count_1_cry_12_TMR_0;
  (* src = "lattice_riscv.v:51067.6-51067.25" *)
  wire main_count_1_cry_12_TMR_1;
  (* src = "lattice_riscv.v:51067.6-51067.25" *)
  wire main_count_1_cry_12_TMR_2;
  (* src = "lattice_riscv.v:50759.6-50759.30" *)
  wire main_count_1_cry_13_0_S0_TMR_0;
  (* src = "lattice_riscv.v:50759.6-50759.30" *)
  wire main_count_1_cry_13_0_S0_TMR_1;
  (* src = "lattice_riscv.v:50759.6-50759.30" *)
  wire main_count_1_cry_13_0_S0_TMR_2;
  (* src = "lattice_riscv.v:50760.6-50760.30" *)
  wire main_count_1_cry_13_0_S1_TMR_0;
  (* src = "lattice_riscv.v:50760.6-50760.30" *)
  wire main_count_1_cry_13_0_S1_TMR_1;
  (* src = "lattice_riscv.v:50760.6-50760.30" *)
  wire main_count_1_cry_13_0_S1_TMR_2;
  (* src = "lattice_riscv.v:51068.6-51068.25" *)
  wire main_count_1_cry_14_TMR_0;
  (* src = "lattice_riscv.v:51068.6-51068.25" *)
  wire main_count_1_cry_14_TMR_1;
  (* src = "lattice_riscv.v:51068.6-51068.25" *)
  wire main_count_1_cry_14_TMR_2;
  (* src = "lattice_riscv.v:50761.6-50761.30" *)
  wire main_count_1_cry_15_0_S0_TMR_0;
  (* src = "lattice_riscv.v:50761.6-50761.30" *)
  wire main_count_1_cry_15_0_S0_TMR_1;
  (* src = "lattice_riscv.v:50761.6-50761.30" *)
  wire main_count_1_cry_15_0_S0_TMR_2;
  (* src = "lattice_riscv.v:50762.6-50762.30" *)
  wire main_count_1_cry_15_0_S1_TMR_0;
  (* src = "lattice_riscv.v:50762.6-50762.30" *)
  wire main_count_1_cry_15_0_S1_TMR_1;
  (* src = "lattice_riscv.v:50762.6-50762.30" *)
  wire main_count_1_cry_15_0_S1_TMR_2;
  (* src = "lattice_riscv.v:51069.6-51069.25" *)
  wire main_count_1_cry_16_TMR_0;
  (* src = "lattice_riscv.v:51069.6-51069.25" *)
  wire main_count_1_cry_16_TMR_1;
  (* src = "lattice_riscv.v:51069.6-51069.25" *)
  wire main_count_1_cry_16_TMR_2;
  (* src = "lattice_riscv.v:50763.6-50763.30" *)
  wire main_count_1_cry_17_0_S0_TMR_0;
  (* src = "lattice_riscv.v:50763.6-50763.30" *)
  wire main_count_1_cry_17_0_S0_TMR_1;
  (* src = "lattice_riscv.v:50763.6-50763.30" *)
  wire main_count_1_cry_17_0_S0_TMR_2;
  (* src = "lattice_riscv.v:50764.6-50764.30" *)
  wire main_count_1_cry_17_0_S1_TMR_0;
  (* src = "lattice_riscv.v:50764.6-50764.30" *)
  wire main_count_1_cry_17_0_S1_TMR_1;
  (* src = "lattice_riscv.v:50764.6-50764.30" *)
  wire main_count_1_cry_17_0_S1_TMR_2;
  (* src = "lattice_riscv.v:51070.6-51070.25" *)
  wire main_count_1_cry_18_TMR_0;
  (* src = "lattice_riscv.v:51070.6-51070.25" *)
  wire main_count_1_cry_18_TMR_1;
  (* src = "lattice_riscv.v:51070.6-51070.25" *)
  wire main_count_1_cry_18_TMR_2;
  (* src = "lattice_riscv.v:50765.6-50765.30" *)
  wire main_count_1_cry_19_0_S0_TMR_0;
  (* src = "lattice_riscv.v:50765.6-50765.30" *)
  wire main_count_1_cry_19_0_S0_TMR_1;
  (* src = "lattice_riscv.v:50765.6-50765.30" *)
  wire main_count_1_cry_19_0_S0_TMR_2;
  (* src = "lattice_riscv.v:50766.6-50766.30" *)
  wire main_count_1_cry_19_0_S1_TMR_0;
  (* src = "lattice_riscv.v:50766.6-50766.30" *)
  wire main_count_1_cry_19_0_S1_TMR_1;
  (* src = "lattice_riscv.v:50766.6-50766.30" *)
  wire main_count_1_cry_19_0_S1_TMR_2;
  (* src = "lattice_riscv.v:50747.6-50747.29" *)
  wire main_count_1_cry_1_0_S0_TMR_0;
  (* src = "lattice_riscv.v:50747.6-50747.29" *)
  wire main_count_1_cry_1_0_S0_TMR_1;
  (* src = "lattice_riscv.v:50747.6-50747.29" *)
  wire main_count_1_cry_1_0_S0_TMR_2;
  (* src = "lattice_riscv.v:50748.6-50748.29" *)
  wire main_count_1_cry_1_0_S1_TMR_0;
  (* src = "lattice_riscv.v:50748.6-50748.29" *)
  wire main_count_1_cry_1_0_S1_TMR_1;
  (* src = "lattice_riscv.v:50748.6-50748.29" *)
  wire main_count_1_cry_1_0_S1_TMR_2;
  (* src = "lattice_riscv.v:51071.6-51071.25" *)
  wire main_count_1_cry_20_TMR_0;
  (* src = "lattice_riscv.v:51071.6-51071.25" *)
  wire main_count_1_cry_20_TMR_1;
  (* src = "lattice_riscv.v:51071.6-51071.25" *)
  wire main_count_1_cry_20_TMR_2;
  (* src = "lattice_riscv.v:51062.6-51062.24" *)
  wire main_count_1_cry_2_TMR_0;
  (* src = "lattice_riscv.v:51062.6-51062.24" *)
  wire main_count_1_cry_2_TMR_1;
  (* src = "lattice_riscv.v:51062.6-51062.24" *)
  wire main_count_1_cry_2_TMR_2;
  (* src = "lattice_riscv.v:50749.6-50749.29" *)
  wire main_count_1_cry_3_0_S0_TMR_0;
  (* src = "lattice_riscv.v:50749.6-50749.29" *)
  wire main_count_1_cry_3_0_S0_TMR_1;
  (* src = "lattice_riscv.v:50749.6-50749.29" *)
  wire main_count_1_cry_3_0_S0_TMR_2;
  (* src = "lattice_riscv.v:50750.6-50750.29" *)
  wire main_count_1_cry_3_0_S1_TMR_0;
  (* src = "lattice_riscv.v:50750.6-50750.29" *)
  wire main_count_1_cry_3_0_S1_TMR_1;
  (* src = "lattice_riscv.v:50750.6-50750.29" *)
  wire main_count_1_cry_3_0_S1_TMR_2;
  (* src = "lattice_riscv.v:51063.6-51063.24" *)
  wire main_count_1_cry_4_TMR_0;
  (* src = "lattice_riscv.v:51063.6-51063.24" *)
  wire main_count_1_cry_4_TMR_1;
  (* src = "lattice_riscv.v:51063.6-51063.24" *)
  wire main_count_1_cry_4_TMR_2;
  (* src = "lattice_riscv.v:50751.6-50751.29" *)
  wire main_count_1_cry_5_0_S0_TMR_0;
  (* src = "lattice_riscv.v:50751.6-50751.29" *)
  wire main_count_1_cry_5_0_S0_TMR_1;
  (* src = "lattice_riscv.v:50751.6-50751.29" *)
  wire main_count_1_cry_5_0_S0_TMR_2;
  (* src = "lattice_riscv.v:50752.6-50752.29" *)
  wire main_count_1_cry_5_0_S1_TMR_0;
  (* src = "lattice_riscv.v:50752.6-50752.29" *)
  wire main_count_1_cry_5_0_S1_TMR_1;
  (* src = "lattice_riscv.v:50752.6-50752.29" *)
  wire main_count_1_cry_5_0_S1_TMR_2;
  (* src = "lattice_riscv.v:51064.6-51064.24" *)
  wire main_count_1_cry_6_TMR_0;
  (* src = "lattice_riscv.v:51064.6-51064.24" *)
  wire main_count_1_cry_6_TMR_1;
  (* src = "lattice_riscv.v:51064.6-51064.24" *)
  wire main_count_1_cry_6_TMR_2;
  (* src = "lattice_riscv.v:50753.6-50753.29" *)
  wire main_count_1_cry_7_0_S0_TMR_0;
  (* src = "lattice_riscv.v:50753.6-50753.29" *)
  wire main_count_1_cry_7_0_S0_TMR_1;
  (* src = "lattice_riscv.v:50753.6-50753.29" *)
  wire main_count_1_cry_7_0_S0_TMR_2;
  (* src = "lattice_riscv.v:50754.6-50754.29" *)
  wire main_count_1_cry_7_0_S1_TMR_0;
  (* src = "lattice_riscv.v:50754.6-50754.29" *)
  wire main_count_1_cry_7_0_S1_TMR_1;
  (* src = "lattice_riscv.v:50754.6-50754.29" *)
  wire main_count_1_cry_7_0_S1_TMR_2;
  (* src = "lattice_riscv.v:51065.6-51065.24" *)
  wire main_count_1_cry_8_TMR_0;
  (* src = "lattice_riscv.v:51065.6-51065.24" *)
  wire main_count_1_cry_8_TMR_1;
  (* src = "lattice_riscv.v:51065.6-51065.24" *)
  wire main_count_1_cry_8_TMR_2;
  (* src = "lattice_riscv.v:50755.6-50755.29" *)
  wire main_count_1_cry_9_0_S0_TMR_0;
  (* src = "lattice_riscv.v:50755.6-50755.29" *)
  wire main_count_1_cry_9_0_S0_TMR_1;
  (* src = "lattice_riscv.v:50755.6-50755.29" *)
  wire main_count_1_cry_9_0_S0_TMR_2;
  (* src = "lattice_riscv.v:50756.6-50756.29" *)
  wire main_count_1_cry_9_0_S1_TMR_0;
  (* src = "lattice_riscv.v:50756.6-50756.29" *)
  wire main_count_1_cry_9_0_S1_TMR_1;
  (* src = "lattice_riscv.v:50756.6-50756.29" *)
  wire main_count_1_cry_9_0_S1_TMR_2;
  (* src = "lattice_riscv.v:51156.6-51156.30" *)
  wire main_count_1_s_21_0_COUT_TMR_0;
  (* src = "lattice_riscv.v:51156.6-51156.30" *)
  wire main_count_1_s_21_0_COUT_TMR_1;
  (* src = "lattice_riscv.v:51156.6-51156.30" *)
  wire main_count_1_s_21_0_COUT_TMR_2;
  (* src = "lattice_riscv.v:50767.6-50767.28" *)
  wire main_count_1_s_21_0_S0_TMR_0;
  (* src = "lattice_riscv.v:50767.6-50767.28" *)
  wire main_count_1_s_21_0_S0_TMR_1;
  (* src = "lattice_riscv.v:50767.6-50767.28" *)
  wire main_count_1_s_21_0_S0_TMR_2;
  (* src = "lattice_riscv.v:51155.6-51155.28" *)
  wire main_count_1_s_21_0_S1_TMR_0;
  (* src = "lattice_riscv.v:51155.6-51155.28" *)
  wire main_count_1_s_21_0_S1_TMR_1;
  (* src = "lattice_riscv.v:51155.6-51155.28" *)
  wire main_count_1_s_21_0_S1_TMR_2;
  (* src = "lattice_riscv.v:50619.13-50619.26" *)
  wire [21:0] main_count_QN;
  (* src = "lattice_riscv.v:50544.12-50544.26" *)
  wire [1:0] main_count_RNO_TMR_0;
  (* src = "lattice_riscv.v:50544.12-50544.26" *)
  wire [1:0] main_count_RNO_TMR_1;
  (* src = "lattice_riscv.v:50544.12-50544.26" *)
  wire [1:0] main_count_RNO_TMR_2;
  (* src = "lattice_riscv.v:50492.13-50492.23" *)
  wire [21:1] main_count_TMR_0;
  (* src = "lattice_riscv.v:50492.13-50492.23" *)
  wire [21:1] main_count_TMR_1;
  (* src = "lattice_riscv.v:50492.13-50492.23" *)
  wire [21:1] main_count_TMR_2;
  (* src = "lattice_riscv.v:50627.14-50627.26" *)
  wire main_count_i_TMR_0;
  (* src = "lattice_riscv.v:50627.14-50627.26" *)
  wire main_count_i_TMR_1;
  (* src = "lattice_riscv.v:50627.14-50627.26" *)
  wire main_count_i_TMR_2;
  (* src = "lattice_riscv.v:50530.13-50530.30" *)
  wire [20:2] main_count_r_0_a2_TMR_0;
  (* src = "lattice_riscv.v:50530.13-50530.30" *)
  wire [20:2] main_count_r_0_a2_TMR_1;
  (* src = "lattice_riscv.v:50530.13-50530.30" *)
  wire [20:2] main_count_r_0_a2_TMR_2;
  (* src = "lattice_riscv.v:50656.6-50656.21" *)
  wire main_crg_clkout;
  (* src = "lattice_riscv.v:50658.6-50658.21" *)
  wire main_crg_locked;
  (* src = "lattice_riscv.v:50620.13-50620.34" *)
  wire [15:0] main_crg_por_count_QN;
  (* src = "lattice_riscv.v:50545.13-50545.35" *)
  wire [15:0] main_crg_por_count_RNO_TMR_0;
  (* src = "lattice_riscv.v:50545.13-50545.35" *)
  wire [15:0] main_crg_por_count_RNO_TMR_1;
  (* src = "lattice_riscv.v:50545.13-50545.35" *)
  wire [15:0] main_crg_por_count_RNO_TMR_2;
  (* src = "lattice_riscv.v:50555.13-50555.31" *)
  wire [15:0] main_crg_por_count_TMR_0;
  (* src = "lattice_riscv.v:50555.13-50555.31" *)
  wire [15:0] main_crg_por_count_TMR_1;
  (* src = "lattice_riscv.v:50555.13-50555.31" *)
  wire [15:0] main_crg_por_count_TMR_2;
  (* src = "lattice_riscv.v:51133.6-51133.26" *)
  wire main_crg_por_done_11_TMR_0;
  (* src = "lattice_riscv.v:51133.6-51133.26" *)
  wire main_crg_por_done_11_TMR_1;
  (* src = "lattice_riscv.v:51133.6-51133.26" *)
  wire main_crg_por_done_11_TMR_2;
  (* src = "lattice_riscv.v:51134.6-51134.26" *)
  wire main_crg_por_done_12_TMR_0;
  (* src = "lattice_riscv.v:51134.6-51134.26" *)
  wire main_crg_por_done_12_TMR_1;
  (* src = "lattice_riscv.v:51134.6-51134.26" *)
  wire main_crg_por_done_12_TMR_2;
  (* src = "lattice_riscv.v:51135.6-51135.26" *)
  wire main_crg_por_done_13_TMR_0;
  (* src = "lattice_riscv.v:51135.6-51135.26" *)
  wire main_crg_por_done_13_TMR_1;
  (* src = "lattice_riscv.v:51135.6-51135.26" *)
  wire main_crg_por_done_13_TMR_2;
  (* src = "lattice_riscv.v:51130.6-51130.25" *)
  wire main_crg_por_done_1_TMR_0;
  (* src = "lattice_riscv.v:51130.6-51130.25" *)
  wire main_crg_por_done_1_TMR_1;
  (* src = "lattice_riscv.v:51130.6-51130.25" *)
  wire main_crg_por_done_1_TMR_2;
  (* src = "lattice_riscv.v:51131.6-51131.25" *)
  wire main_crg_por_done_5_TMR_0;
  (* src = "lattice_riscv.v:51131.6-51131.25" *)
  wire main_crg_por_done_5_TMR_1;
  (* src = "lattice_riscv.v:51131.6-51131.25" *)
  wire main_crg_por_done_5_TMR_2;
  (* src = "lattice_riscv.v:51132.6-51132.25" *)
  wire main_crg_por_done_9_TMR_0;
  (* src = "lattice_riscv.v:51132.6-51132.25" *)
  wire main_crg_por_done_9_TMR_1;
  (* src = "lattice_riscv.v:51132.6-51132.25" *)
  wire main_crg_por_done_9_TMR_2;
  wire main_cs06_0_RED_VOTER_wire;
  (* src = "lattice_riscv.v:50731.6-50731.15" *)
  wire main_cs06_TMR_0;
  (* src = "lattice_riscv.v:50731.6-50731.15" *)
  wire main_cs06_TMR_1;
  (* src = "lattice_riscv.v:50731.6-50731.15" *)
  wire main_cs06_TMR_2;
  (* src = "lattice_riscv.v:50488.13-50488.26" *)
  wire [31:0] main_dataout0;
  (* src = "lattice_riscv.v:50489.13-50489.26" *)
  wire [31:0] main_dataout1;
  (* src = "lattice_riscv.v:51137.6-51137.18" *)
  wire main_done_11_TMR_0;
  (* src = "lattice_riscv.v:51137.6-51137.18" *)
  wire main_done_11_TMR_1;
  (* src = "lattice_riscv.v:51137.6-51137.18" *)
  wire main_done_11_TMR_2;
  (* src = "lattice_riscv.v:51138.6-51138.18" *)
  wire main_done_12_TMR_0;
  (* src = "lattice_riscv.v:51138.6-51138.18" *)
  wire main_done_12_TMR_1;
  (* src = "lattice_riscv.v:51138.6-51138.18" *)
  wire main_done_12_TMR_2;
  (* src = "lattice_riscv.v:51139.6-51139.18" *)
  wire main_done_13_TMR_0;
  (* src = "lattice_riscv.v:51139.6-51139.18" *)
  wire main_done_13_TMR_1;
  (* src = "lattice_riscv.v:51139.6-51139.18" *)
  wire main_done_13_TMR_2;
  (* src = "lattice_riscv.v:51140.6-51140.18" *)
  wire main_done_15_TMR_0;
  (* src = "lattice_riscv.v:51140.6-51140.18" *)
  wire main_done_15_TMR_1;
  (* src = "lattice_riscv.v:51140.6-51140.18" *)
  wire main_done_15_TMR_2;
  (* src = "lattice_riscv.v:51141.6-51141.18" *)
  wire main_done_16_TMR_0;
  (* src = "lattice_riscv.v:51141.6-51141.18" *)
  wire main_done_16_TMR_1;
  (* src = "lattice_riscv.v:51141.6-51141.18" *)
  wire main_done_16_TMR_2;
  (* src = "lattice_riscv.v:51142.6-51142.18" *)
  wire main_done_18_TMR_0;
  (* src = "lattice_riscv.v:51142.6-51142.18" *)
  wire main_done_18_TMR_1;
  (* src = "lattice_riscv.v:51142.6-51142.18" *)
  wire main_done_18_TMR_2;
  (* src = "lattice_riscv.v:51136.6-51136.17" *)
  wire main_done_7_TMR_0;
  (* src = "lattice_riscv.v:51136.6-51136.17" *)
  wire main_done_7_TMR_1;
  (* src = "lattice_riscv.v:51136.6-51136.17" *)
  wire main_done_7_TMR_2;
  (* src = "lattice_riscv.v:50695.6-50695.15" *)
  wire main_done_TMR_0;
  (* src = "lattice_riscv.v:50695.6-50695.15" *)
  wire main_done_TMR_1;
  (* src = "lattice_riscv.v:50695.6-50695.15" *)
  wire main_done_TMR_2;
  (* src = "lattice_riscv.v:51246.6-51246.21" *)
  wire \main_mode.fb_0_TMR_0 ;
  (* src = "lattice_riscv.v:51246.6-51246.21" *)
  wire \main_mode.fb_0_TMR_1 ;
  (* src = "lattice_riscv.v:51246.6-51246.21" *)
  wire \main_mode.fb_0_TMR_2 ;
  (* src = "lattice_riscv.v:51232.6-51232.18" *)
  wire main_mode_QN;
  (* src = "lattice_riscv.v:50686.6-50686.15" *)
  wire main_mode_TMR_0;
  (* src = "lattice_riscv.v:50686.6-50686.15" *)
  wire main_mode_TMR_1;
  (* src = "lattice_riscv.v:50686.6-50686.15" *)
  wire main_mode_TMR_2;
  (* src = "lattice_riscv.v:51233.6-51233.16" *)
  wire main_re_QN;
  (* src = "lattice_riscv.v:50720.6-50720.13" *)
  wire main_re_TMR_0;
  (* src = "lattice_riscv.v:50720.6-50720.13" *)
  wire main_re_TMR_1;
  (* src = "lattice_riscv.v:50720.6-50720.13" *)
  wire main_re_TMR_2;
  (* src = "lattice_riscv.v:50714.6-50714.27" *)
  wire main_storage_0_sqmuxa_TMR_0;
  (* src = "lattice_riscv.v:50714.6-50714.27" *)
  wire main_storage_0_sqmuxa_TMR_1;
  (* src = "lattice_riscv.v:50714.6-50714.27" *)
  wire main_storage_0_sqmuxa_TMR_2;
  (* src = "lattice_riscv.v:50621.13-50621.28" *)
  wire [13:0] main_storage_QN;
  (* src = "lattice_riscv.v:50498.13-50498.25" *)
  wire [13:0] main_storage_TMR_0;
  (* src = "lattice_riscv.v:50498.13-50498.25" *)
  wire [13:0] main_storage_TMR_1;
  (* src = "lattice_riscv.v:50498.13-50498.25" *)
  wire [13:0] main_storage_TMR_2;
  wire main_wren0_0_RED_VOTER_wire;
  (* src = "lattice_riscv.v:50654.6-50654.16" *)
  wire main_wren0_TMR_0;
  (* src = "lattice_riscv.v:50654.6-50654.16" *)
  wire main_wren0_TMR_1;
  (* src = "lattice_riscv.v:50654.6-50654.16" *)
  wire main_wren0_TMR_2;
  wire main_wren1_0_RED_VOTER_wire;
  (* src = "lattice_riscv.v:50655.6-50655.16" *)
  wire main_wren1_TMR_0;
  (* src = "lattice_riscv.v:50655.6-50655.16" *)
  wire main_wren1_TMR_1;
  (* src = "lattice_riscv.v:50655.6-50655.16" *)
  wire main_wren1_TMR_2;
  (* src = "lattice_riscv.v:50622.12-50622.23" *)
  wire [5:0] mem_adr0_QN;
  (* src = "lattice_riscv.v:50495.12-50495.20" *)
  wire [5:0] mem_adr0_TMR_0;
  (* src = "lattice_riscv.v:50495.12-50495.20" *)
  wire [5:0] mem_adr0_TMR_1;
  (* src = "lattice_riscv.v:50495.12-50495.20" *)
  wire [5:0] mem_adr0_TMR_2;
  (* src = "lattice_riscv.v:50660.6-50660.13" *)
  wire por_rst_TMR_0;
  (* src = "lattice_riscv.v:50660.6-50660.13" *)
  wire por_rst_TMR_1;
  (* src = "lattice_riscv.v:50660.6-50660.13" *)
  wire por_rst_TMR_2;
  (* src = "lattice_riscv.v:50501.13-50501.21" *)
  wire [31:0] rom_dat0;
  (* src = "lattice_riscv.v:50565.13-50565.30" *)
  wire [17:2] rom_dat0_2_0_0_DO;
  (* src = "lattice_riscv.v:50575.13-50575.31" *)
  wire [17:2] rom_dat0_2_0_10_DO;
  (* src = "lattice_riscv.v:50576.13-50576.31" *)
  wire [17:2] rom_dat0_2_0_11_DO;
  (* src = "lattice_riscv.v:50577.13-50577.31" *)
  wire [17:2] rom_dat0_2_0_12_DO;
  (* src = "lattice_riscv.v:50578.13-50578.31" *)
  wire [17:2] rom_dat0_2_0_13_DO;
  (* src = "lattice_riscv.v:50579.13-50579.31" *)
  wire [17:2] rom_dat0_2_0_14_DO;
  (* src = "lattice_riscv.v:50580.13-50580.31" *)
  wire [17:2] rom_dat0_2_0_15_DO;
  (* src = "lattice_riscv.v:50566.13-50566.30" *)
  wire [17:2] rom_dat0_2_0_1_DO;
  (* src = "lattice_riscv.v:50567.13-50567.30" *)
  wire [17:2] rom_dat0_2_0_2_DO;
  (* src = "lattice_riscv.v:50568.13-50568.30" *)
  wire [17:2] rom_dat0_2_0_3_DO;
  (* src = "lattice_riscv.v:50569.13-50569.30" *)
  wire [17:2] rom_dat0_2_0_4_DO;
  (* src = "lattice_riscv.v:50570.13-50570.30" *)
  wire [17:2] rom_dat0_2_0_5_DO;
  (* src = "lattice_riscv.v:50571.13-50571.30" *)
  wire [17:2] rom_dat0_2_0_6_DO;
  (* src = "lattice_riscv.v:50572.13-50572.30" *)
  wire [17:2] rom_dat0_2_0_7_DO;
  (* src = "lattice_riscv.v:50573.13-50573.30" *)
  wire [17:2] rom_dat0_2_0_8_DO;
  (* src = "lattice_riscv.v:50574.13-50574.30" *)
  wire [17:2] rom_dat0_2_0_9_DO;
  (* src = "lattice_riscv.v:50448.7-50448.16" *)
  input serial_rx;
  wire serial_rx;
  (* src = "lattice_riscv.v:51186.6-51186.17" *)
  wire serial_rx_c;
  (* src = "lattice_riscv.v:50449.8-50449.17" *)
  output serial_tx;
  wire serial_tx;
  (* src = "lattice_riscv.v:50697.6-50697.17" *)
  wire serial_tx_4_TMR_0;
  (* src = "lattice_riscv.v:50697.6-50697.17" *)
  wire serial_tx_4_TMR_1;
  (* src = "lattice_riscv.v:50697.6-50697.17" *)
  wire serial_tx_4_TMR_2;
  wire serial_tx_c_0_RED_VOTER_wire;
  (* src = "lattice_riscv.v:51187.6-51187.17" *)
  wire serial_tx_c_TMR_0;
  (* src = "lattice_riscv.v:51187.6-51187.17" *)
  wire serial_tx_c_TMR_1;
  (* src = "lattice_riscv.v:51187.6-51187.17" *)
  wire serial_tx_c_TMR_2;
  (* src = "lattice_riscv.v:50512.12-50512.21" *)
  wire [7:0] storage_1_TMR_0;
  (* src = "lattice_riscv.v:50512.12-50512.21" *)
  wire [7:0] storage_1_TMR_1;
  (* src = "lattice_riscv.v:50512.12-50512.21" *)
  wire [7:0] storage_1_TMR_2;
  (* src = "lattice_riscv.v:50623.12-50623.29" *)
  wire [7:0] storage_1_dat1_QN;
  (* src = "lattice_riscv.v:50515.12-50515.26" *)
  wire [7:0] storage_1_dat1_TMR_0;
  (* src = "lattice_riscv.v:50515.12-50515.26" *)
  wire [7:0] storage_1_dat1_TMR_1;
  (* src = "lattice_riscv.v:50515.12-50515.26" *)
  wire [7:0] storage_1_dat1_TMR_2;
  (* src = "lattice_riscv.v:50523.12-50523.19" *)
  wire [7:0] storage_TMR_0;
  (* src = "lattice_riscv.v:50523.12-50523.19" *)
  wire [7:0] storage_TMR_1;
  (* src = "lattice_riscv.v:50523.12-50523.19" *)
  wire [7:0] storage_TMR_2;
  (* src = "lattice_riscv.v:50624.12-50624.27" *)
  wire [7:0] storage_dat1_QN;
  (* src = "lattice_riscv.v:50506.12-50506.24" *)
  wire [7:0] storage_dat1_TMR_0;
  (* src = "lattice_riscv.v:50506.12-50506.24" *)
  wire [7:0] storage_dat1_TMR_1;
  (* src = "lattice_riscv.v:50506.12-50506.24" *)
  wire [7:0] storage_dat1_TMR_2;
  (* src = "lattice_riscv.v:50487.12-50487.19" *)
  wire sys_clk;
  (* src = "lattice_riscv.v:50662.6-50662.13" *)
  wire sys_rst_TMR_0;
  (* src = "lattice_riscv.v:50662.6-50662.13" *)
  wire sys_rst_TMR_1;
  (* src = "lattice_riscv.v:50662.6-50662.13" *)
  wire sys_rst_TMR_2;
  (* src = "lattice_riscv.v:50537.13-50537.44" *)
  wire [31:0] un1_main_basesoc_bus_errors_1_0_TMR_0;
  (* src = "lattice_riscv.v:50537.13-50537.44" *)
  wire [31:0] un1_main_basesoc_bus_errors_1_0_TMR_1;
  (* src = "lattice_riscv.v:50537.13-50537.44" *)
  wire [31:0] un1_main_basesoc_bus_errors_1_0_TMR_2;
  (* src = "lattice_riscv.v:50558.13-50558.42" *)
  wire [31:0] un1_main_basesoc_bus_errors_1_TMR_0;
  (* src = "lattice_riscv.v:50558.13-50558.42" *)
  wire [31:0] un1_main_basesoc_bus_errors_1_TMR_1;
  (* src = "lattice_riscv.v:50558.13-50558.42" *)
  wire [31:0] un1_main_basesoc_bus_errors_1_TMR_2;
  (* src = "lattice_riscv.v:51167.6-51167.46" *)
  wire un1_main_basesoc_bus_errors_1_cry_0_0_S0_TMR_0;
  (* src = "lattice_riscv.v:51167.6-51167.46" *)
  wire un1_main_basesoc_bus_errors_1_cry_0_0_S0_TMR_1;
  (* src = "lattice_riscv.v:51167.6-51167.46" *)
  wire un1_main_basesoc_bus_errors_1_cry_0_0_S0_TMR_2;
  (* src = "lattice_riscv.v:50995.6-50995.41" *)
  wire un1_main_basesoc_bus_errors_1_cry_0_TMR_0;
  (* src = "lattice_riscv.v:50995.6-50995.41" *)
  wire un1_main_basesoc_bus_errors_1_cry_0_TMR_1;
  (* src = "lattice_riscv.v:50995.6-50995.41" *)
  wire un1_main_basesoc_bus_errors_1_cry_0_TMR_2;
  (* src = "lattice_riscv.v:51000.6-51000.42" *)
  wire un1_main_basesoc_bus_errors_1_cry_10_TMR_0;
  (* src = "lattice_riscv.v:51000.6-51000.42" *)
  wire un1_main_basesoc_bus_errors_1_cry_10_TMR_1;
  (* src = "lattice_riscv.v:51000.6-51000.42" *)
  wire un1_main_basesoc_bus_errors_1_cry_10_TMR_2;
  (* src = "lattice_riscv.v:51001.6-51001.42" *)
  wire un1_main_basesoc_bus_errors_1_cry_12_TMR_0;
  (* src = "lattice_riscv.v:51001.6-51001.42" *)
  wire un1_main_basesoc_bus_errors_1_cry_12_TMR_1;
  (* src = "lattice_riscv.v:51001.6-51001.42" *)
  wire un1_main_basesoc_bus_errors_1_cry_12_TMR_2;
  (* src = "lattice_riscv.v:51002.6-51002.42" *)
  wire un1_main_basesoc_bus_errors_1_cry_14_TMR_0;
  (* src = "lattice_riscv.v:51002.6-51002.42" *)
  wire un1_main_basesoc_bus_errors_1_cry_14_TMR_1;
  (* src = "lattice_riscv.v:51002.6-51002.42" *)
  wire un1_main_basesoc_bus_errors_1_cry_14_TMR_2;
  (* src = "lattice_riscv.v:51003.6-51003.42" *)
  wire un1_main_basesoc_bus_errors_1_cry_16_TMR_0;
  (* src = "lattice_riscv.v:51003.6-51003.42" *)
  wire un1_main_basesoc_bus_errors_1_cry_16_TMR_1;
  (* src = "lattice_riscv.v:51003.6-51003.42" *)
  wire un1_main_basesoc_bus_errors_1_cry_16_TMR_2;
  (* src = "lattice_riscv.v:51004.6-51004.42" *)
  wire un1_main_basesoc_bus_errors_1_cry_18_TMR_0;
  (* src = "lattice_riscv.v:51004.6-51004.42" *)
  wire un1_main_basesoc_bus_errors_1_cry_18_TMR_1;
  (* src = "lattice_riscv.v:51004.6-51004.42" *)
  wire un1_main_basesoc_bus_errors_1_cry_18_TMR_2;
  (* src = "lattice_riscv.v:51005.6-51005.42" *)
  wire un1_main_basesoc_bus_errors_1_cry_20_TMR_0;
  (* src = "lattice_riscv.v:51005.6-51005.42" *)
  wire un1_main_basesoc_bus_errors_1_cry_20_TMR_1;
  (* src = "lattice_riscv.v:51005.6-51005.42" *)
  wire un1_main_basesoc_bus_errors_1_cry_20_TMR_2;
  (* src = "lattice_riscv.v:51006.6-51006.42" *)
  wire un1_main_basesoc_bus_errors_1_cry_22_TMR_0;
  (* src = "lattice_riscv.v:51006.6-51006.42" *)
  wire un1_main_basesoc_bus_errors_1_cry_22_TMR_1;
  (* src = "lattice_riscv.v:51006.6-51006.42" *)
  wire un1_main_basesoc_bus_errors_1_cry_22_TMR_2;
  (* src = "lattice_riscv.v:51007.6-51007.42" *)
  wire un1_main_basesoc_bus_errors_1_cry_24_TMR_0;
  (* src = "lattice_riscv.v:51007.6-51007.42" *)
  wire un1_main_basesoc_bus_errors_1_cry_24_TMR_1;
  (* src = "lattice_riscv.v:51007.6-51007.42" *)
  wire un1_main_basesoc_bus_errors_1_cry_24_TMR_2;
  (* src = "lattice_riscv.v:51008.6-51008.42" *)
  wire un1_main_basesoc_bus_errors_1_cry_26_TMR_0;
  (* src = "lattice_riscv.v:51008.6-51008.42" *)
  wire un1_main_basesoc_bus_errors_1_cry_26_TMR_1;
  (* src = "lattice_riscv.v:51008.6-51008.42" *)
  wire un1_main_basesoc_bus_errors_1_cry_26_TMR_2;
  (* src = "lattice_riscv.v:51009.6-51009.42" *)
  wire un1_main_basesoc_bus_errors_1_cry_28_TMR_0;
  (* src = "lattice_riscv.v:51009.6-51009.42" *)
  wire un1_main_basesoc_bus_errors_1_cry_28_TMR_1;
  (* src = "lattice_riscv.v:51009.6-51009.42" *)
  wire un1_main_basesoc_bus_errors_1_cry_28_TMR_2;
  (* src = "lattice_riscv.v:50996.6-50996.41" *)
  wire un1_main_basesoc_bus_errors_1_cry_2_TMR_0;
  (* src = "lattice_riscv.v:50996.6-50996.41" *)
  wire un1_main_basesoc_bus_errors_1_cry_2_TMR_1;
  (* src = "lattice_riscv.v:50996.6-50996.41" *)
  wire un1_main_basesoc_bus_errors_1_cry_2_TMR_2;
  (* src = "lattice_riscv.v:51010.6-51010.42" *)
  wire un1_main_basesoc_bus_errors_1_cry_30_TMR_0;
  (* src = "lattice_riscv.v:51010.6-51010.42" *)
  wire un1_main_basesoc_bus_errors_1_cry_30_TMR_1;
  (* src = "lattice_riscv.v:51010.6-51010.42" *)
  wire un1_main_basesoc_bus_errors_1_cry_30_TMR_2;
  (* src = "lattice_riscv.v:50997.6-50997.41" *)
  wire un1_main_basesoc_bus_errors_1_cry_4_TMR_0;
  (* src = "lattice_riscv.v:50997.6-50997.41" *)
  wire un1_main_basesoc_bus_errors_1_cry_4_TMR_1;
  (* src = "lattice_riscv.v:50997.6-50997.41" *)
  wire un1_main_basesoc_bus_errors_1_cry_4_TMR_2;
  (* src = "lattice_riscv.v:50998.6-50998.41" *)
  wire un1_main_basesoc_bus_errors_1_cry_6_TMR_0;
  (* src = "lattice_riscv.v:50998.6-50998.41" *)
  wire un1_main_basesoc_bus_errors_1_cry_6_TMR_1;
  (* src = "lattice_riscv.v:50998.6-50998.41" *)
  wire un1_main_basesoc_bus_errors_1_cry_6_TMR_2;
  (* src = "lattice_riscv.v:50999.6-50999.41" *)
  wire un1_main_basesoc_bus_errors_1_cry_8_TMR_0;
  (* src = "lattice_riscv.v:50999.6-50999.41" *)
  wire un1_main_basesoc_bus_errors_1_cry_8_TMR_1;
  (* src = "lattice_riscv.v:50999.6-50999.41" *)
  wire un1_main_basesoc_bus_errors_1_cry_8_TMR_2;
  (* src = "lattice_riscv.v:51169.6-51169.47" *)
  wire un1_main_basesoc_bus_errors_1_s_31_0_COUT_TMR_0;
  (* src = "lattice_riscv.v:51169.6-51169.47" *)
  wire un1_main_basesoc_bus_errors_1_s_31_0_COUT_TMR_1;
  (* src = "lattice_riscv.v:51169.6-51169.47" *)
  wire un1_main_basesoc_bus_errors_1_s_31_0_COUT_TMR_2;
  (* src = "lattice_riscv.v:51168.6-51168.45" *)
  wire un1_main_basesoc_bus_errors_1_s_31_0_S1_TMR_0;
  (* src = "lattice_riscv.v:51168.6-51168.45" *)
  wire un1_main_basesoc_bus_errors_1_s_31_0_S1_TMR_1;
  (* src = "lattice_riscv.v:51168.6-51168.45" *)
  wire un1_main_basesoc_bus_errors_1_s_31_0_S1_TMR_2;
  (* src = "lattice_riscv.v:50564.12-50564.65" *)
  wire un1_main_basesoc_serial_tx_rs232phytx_next_value112_i_TMR_0;
  (* src = "lattice_riscv.v:50564.12-50564.65" *)
  wire un1_main_basesoc_serial_tx_rs232phytx_next_value112_i_TMR_1;
  (* src = "lattice_riscv.v:50564.12-50564.65" *)
  wire un1_main_basesoc_serial_tx_rs232phytx_next_value112_i_TMR_2;
  (* src = "lattice_riscv.v:51072.6-51072.50" *)
  wire un1_main_basesoc_uart_rx_fifo_consume_axbxc0_TMR_0;
  (* src = "lattice_riscv.v:51072.6-51072.50" *)
  wire un1_main_basesoc_uart_rx_fifo_consume_axbxc0_TMR_1;
  (* src = "lattice_riscv.v:51072.6-51072.50" *)
  wire un1_main_basesoc_uart_rx_fifo_consume_axbxc0_TMR_2;
  (* src = "lattice_riscv.v:51073.6-51073.50" *)
  wire un1_main_basesoc_uart_rx_fifo_consume_axbxc1_TMR_0;
  (* src = "lattice_riscv.v:51073.6-51073.50" *)
  wire un1_main_basesoc_uart_rx_fifo_consume_axbxc1_TMR_1;
  (* src = "lattice_riscv.v:51073.6-51073.50" *)
  wire un1_main_basesoc_uart_rx_fifo_consume_axbxc1_TMR_2;
  (* src = "lattice_riscv.v:51074.6-51074.50" *)
  wire un1_main_basesoc_uart_rx_fifo_consume_axbxc3_TMR_0;
  (* src = "lattice_riscv.v:51074.6-51074.50" *)
  wire un1_main_basesoc_uart_rx_fifo_consume_axbxc3_TMR_1;
  (* src = "lattice_riscv.v:51074.6-51074.50" *)
  wire un1_main_basesoc_uart_rx_fifo_consume_axbxc3_TMR_2;
  (* src = "lattice_riscv.v:51075.6-51075.46" *)
  wire un1_main_basesoc_uart_rx_fifo_consume_c2_TMR_0;
  (* src = "lattice_riscv.v:51075.6-51075.46" *)
  wire un1_main_basesoc_uart_rx_fifo_consume_c2_TMR_1;
  (* src = "lattice_riscv.v:51075.6-51075.46" *)
  wire un1_main_basesoc_uart_rx_fifo_consume_c2_TMR_2;
  (* src = "lattice_riscv.v:50540.12-50540.50" *)
  wire [4:1] un1_main_basesoc_uart_rx_fifo_level0_0_TMR_0;
  (* src = "lattice_riscv.v:50540.12-50540.50" *)
  wire [4:1] un1_main_basesoc_uart_rx_fifo_level0_0_TMR_1;
  (* src = "lattice_riscv.v:50540.12-50540.50" *)
  wire [4:1] un1_main_basesoc_uart_rx_fifo_level0_0_TMR_2;
  (* src = "lattice_riscv.v:50541.12-50541.48" *)
  wire [4:1] un1_main_basesoc_uart_rx_fifo_level0_TMR_0;
  (* src = "lattice_riscv.v:50541.12-50541.48" *)
  wire [4:1] un1_main_basesoc_uart_rx_fifo_level0_TMR_1;
  (* src = "lattice_riscv.v:50541.12-50541.48" *)
  wire [4:1] un1_main_basesoc_uart_rx_fifo_level0_TMR_2;
  (* src = "lattice_riscv.v:51173.6-51173.53" *)
  wire un1_main_basesoc_uart_rx_fifo_level0_cry_0_0_S0_TMR_0;
  (* src = "lattice_riscv.v:51173.6-51173.53" *)
  wire un1_main_basesoc_uart_rx_fifo_level0_cry_0_0_S0_TMR_1;
  (* src = "lattice_riscv.v:51173.6-51173.53" *)
  wire un1_main_basesoc_uart_rx_fifo_level0_cry_0_0_S0_TMR_2;
  (* src = "lattice_riscv.v:51153.6-51153.53" *)
  wire un1_main_basesoc_uart_rx_fifo_level0_cry_0_0_S1_TMR_0;
  (* src = "lattice_riscv.v:51153.6-51153.53" *)
  wire un1_main_basesoc_uart_rx_fifo_level0_cry_0_0_S1_TMR_1;
  (* src = "lattice_riscv.v:51153.6-51153.53" *)
  wire un1_main_basesoc_uart_rx_fifo_level0_cry_0_0_S1_TMR_2;
  (* src = "lattice_riscv.v:50991.6-50991.48" *)
  wire un1_main_basesoc_uart_rx_fifo_level0_cry_0_TMR_0;
  (* src = "lattice_riscv.v:50991.6-50991.48" *)
  wire un1_main_basesoc_uart_rx_fifo_level0_cry_0_TMR_1;
  (* src = "lattice_riscv.v:50991.6-50991.48" *)
  wire un1_main_basesoc_uart_rx_fifo_level0_cry_0_TMR_2;
  (* src = "lattice_riscv.v:50992.6-50992.48" *)
  wire un1_main_basesoc_uart_rx_fifo_level0_cry_2_TMR_0;
  (* src = "lattice_riscv.v:50992.6-50992.48" *)
  wire un1_main_basesoc_uart_rx_fifo_level0_cry_2_TMR_1;
  (* src = "lattice_riscv.v:50992.6-50992.48" *)
  wire un1_main_basesoc_uart_rx_fifo_level0_cry_2_TMR_2;
  (* src = "lattice_riscv.v:51174.6-51174.55" *)
  wire un1_main_basesoc_uart_rx_fifo_level0_cry_3_0_COUT_TMR_0;
  (* src = "lattice_riscv.v:51174.6-51174.55" *)
  wire un1_main_basesoc_uart_rx_fifo_level0_cry_3_0_COUT_TMR_1;
  (* src = "lattice_riscv.v:51174.6-51174.55" *)
  wire un1_main_basesoc_uart_rx_fifo_level0_cry_3_0_COUT_TMR_2;
  (* src = "lattice_riscv.v:50988.6-50988.49" *)
  wire un1_main_basesoc_uart_rx_fifo_level0_scalar_TMR_0;
  (* src = "lattice_riscv.v:50988.6-50988.49" *)
  wire un1_main_basesoc_uart_rx_fifo_level0_scalar_TMR_1;
  (* src = "lattice_riscv.v:50988.6-50988.49" *)
  wire un1_main_basesoc_uart_rx_fifo_level0_scalar_TMR_2;
  (* src = "lattice_riscv.v:51080.6-51080.50" *)
  wire un1_main_basesoc_uart_rx_fifo_produce_axbxc0_TMR_0;
  (* src = "lattice_riscv.v:51080.6-51080.50" *)
  wire un1_main_basesoc_uart_rx_fifo_produce_axbxc0_TMR_1;
  (* src = "lattice_riscv.v:51080.6-51080.50" *)
  wire un1_main_basesoc_uart_rx_fifo_produce_axbxc0_TMR_2;
  (* src = "lattice_riscv.v:51081.6-51081.50" *)
  wire un1_main_basesoc_uart_rx_fifo_produce_axbxc1_TMR_0;
  (* src = "lattice_riscv.v:51081.6-51081.50" *)
  wire un1_main_basesoc_uart_rx_fifo_produce_axbxc1_TMR_1;
  (* src = "lattice_riscv.v:51081.6-51081.50" *)
  wire un1_main_basesoc_uart_rx_fifo_produce_axbxc1_TMR_2;
  (* src = "lattice_riscv.v:51082.6-51082.50" *)
  wire un1_main_basesoc_uart_rx_fifo_produce_axbxc3_TMR_0;
  (* src = "lattice_riscv.v:51082.6-51082.50" *)
  wire un1_main_basesoc_uart_rx_fifo_produce_axbxc3_TMR_1;
  (* src = "lattice_riscv.v:51082.6-51082.50" *)
  wire un1_main_basesoc_uart_rx_fifo_produce_axbxc3_TMR_2;
  (* src = "lattice_riscv.v:51083.6-51083.46" *)
  wire un1_main_basesoc_uart_rx_fifo_produce_c2_TMR_0;
  (* src = "lattice_riscv.v:51083.6-51083.46" *)
  wire un1_main_basesoc_uart_rx_fifo_produce_c2_TMR_1;
  (* src = "lattice_riscv.v:51083.6-51083.46" *)
  wire un1_main_basesoc_uart_rx_fifo_produce_c2_TMR_2;
  (* src = "lattice_riscv.v:51076.6-51076.50" *)
  wire un1_main_basesoc_uart_tx_fifo_consume_axbxc0_TMR_0;
  (* src = "lattice_riscv.v:51076.6-51076.50" *)
  wire un1_main_basesoc_uart_tx_fifo_consume_axbxc0_TMR_1;
  (* src = "lattice_riscv.v:51076.6-51076.50" *)
  wire un1_main_basesoc_uart_tx_fifo_consume_axbxc0_TMR_2;
  (* src = "lattice_riscv.v:51077.6-51077.50" *)
  wire un1_main_basesoc_uart_tx_fifo_consume_axbxc1_TMR_0;
  (* src = "lattice_riscv.v:51077.6-51077.50" *)
  wire un1_main_basesoc_uart_tx_fifo_consume_axbxc1_TMR_1;
  (* src = "lattice_riscv.v:51077.6-51077.50" *)
  wire un1_main_basesoc_uart_tx_fifo_consume_axbxc1_TMR_2;
  (* src = "lattice_riscv.v:51078.6-51078.50" *)
  wire un1_main_basesoc_uart_tx_fifo_consume_axbxc3_TMR_0;
  (* src = "lattice_riscv.v:51078.6-51078.50" *)
  wire un1_main_basesoc_uart_tx_fifo_consume_axbxc3_TMR_1;
  (* src = "lattice_riscv.v:51078.6-51078.50" *)
  wire un1_main_basesoc_uart_tx_fifo_consume_axbxc3_TMR_2;
  (* src = "lattice_riscv.v:51079.6-51079.46" *)
  wire un1_main_basesoc_uart_tx_fifo_consume_c2_TMR_0;
  (* src = "lattice_riscv.v:51079.6-51079.46" *)
  wire un1_main_basesoc_uart_tx_fifo_consume_c2_TMR_1;
  (* src = "lattice_riscv.v:51079.6-51079.46" *)
  wire un1_main_basesoc_uart_tx_fifo_consume_c2_TMR_2;
  (* src = "lattice_riscv.v:50542.12-50542.50" *)
  wire [4:1] un1_main_basesoc_uart_tx_fifo_level0_0_TMR_0;
  (* src = "lattice_riscv.v:50542.12-50542.50" *)
  wire [4:1] un1_main_basesoc_uart_tx_fifo_level0_0_TMR_1;
  (* src = "lattice_riscv.v:50542.12-50542.50" *)
  wire [4:1] un1_main_basesoc_uart_tx_fifo_level0_0_TMR_2;
  (* src = "lattice_riscv.v:50543.12-50543.48" *)
  wire [4:0] un1_main_basesoc_uart_tx_fifo_level0_TMR_0;
  (* src = "lattice_riscv.v:50543.12-50543.48" *)
  wire [4:0] un1_main_basesoc_uart_tx_fifo_level0_TMR_1;
  (* src = "lattice_riscv.v:50543.12-50543.48" *)
  wire [4:0] un1_main_basesoc_uart_tx_fifo_level0_TMR_2;
  (* src = "lattice_riscv.v:51170.6-51170.53" *)
  wire un1_main_basesoc_uart_tx_fifo_level0_cry_0_0_S0_TMR_0;
  (* src = "lattice_riscv.v:51170.6-51170.53" *)
  wire un1_main_basesoc_uart_tx_fifo_level0_cry_0_0_S0_TMR_1;
  (* src = "lattice_riscv.v:51170.6-51170.53" *)
  wire un1_main_basesoc_uart_tx_fifo_level0_cry_0_0_S0_TMR_2;
  (* src = "lattice_riscv.v:51171.6-51171.53" *)
  wire un1_main_basesoc_uart_tx_fifo_level0_cry_0_0_S1_TMR_0;
  (* src = "lattice_riscv.v:51171.6-51171.53" *)
  wire un1_main_basesoc_uart_tx_fifo_level0_cry_0_0_S1_TMR_1;
  (* src = "lattice_riscv.v:51171.6-51171.53" *)
  wire un1_main_basesoc_uart_tx_fifo_level0_cry_0_0_S1_TMR_2;
  (* src = "lattice_riscv.v:50993.6-50993.48" *)
  wire un1_main_basesoc_uart_tx_fifo_level0_cry_0_TMR_0;
  (* src = "lattice_riscv.v:50993.6-50993.48" *)
  wire un1_main_basesoc_uart_tx_fifo_level0_cry_0_TMR_1;
  (* src = "lattice_riscv.v:50993.6-50993.48" *)
  wire un1_main_basesoc_uart_tx_fifo_level0_cry_0_TMR_2;
  (* src = "lattice_riscv.v:50994.6-50994.48" *)
  wire un1_main_basesoc_uart_tx_fifo_level0_cry_2_TMR_0;
  (* src = "lattice_riscv.v:50994.6-50994.48" *)
  wire un1_main_basesoc_uart_tx_fifo_level0_cry_2_TMR_1;
  (* src = "lattice_riscv.v:50994.6-50994.48" *)
  wire un1_main_basesoc_uart_tx_fifo_level0_cry_2_TMR_2;
  (* src = "lattice_riscv.v:51172.6-51172.55" *)
  wire un1_main_basesoc_uart_tx_fifo_level0_cry_3_0_COUT_TMR_0;
  (* src = "lattice_riscv.v:51172.6-51172.55" *)
  wire un1_main_basesoc_uart_tx_fifo_level0_cry_3_0_COUT_TMR_1;
  (* src = "lattice_riscv.v:51172.6-51172.55" *)
  wire un1_main_basesoc_uart_tx_fifo_level0_cry_3_0_COUT_TMR_2;
  (* src = "lattice_riscv.v:50987.6-50987.49" *)
  wire un1_main_basesoc_uart_tx_fifo_level0_scalar_TMR_0;
  (* src = "lattice_riscv.v:50987.6-50987.49" *)
  wire un1_main_basesoc_uart_tx_fifo_level0_scalar_TMR_1;
  (* src = "lattice_riscv.v:50987.6-50987.49" *)
  wire un1_main_basesoc_uart_tx_fifo_level0_scalar_TMR_2;
  (* src = "lattice_riscv.v:51147.6-51147.49" *)
  wire un1_main_basesoc_uart_tx_fifo_produce_ac0_0_TMR_0;
  (* src = "lattice_riscv.v:51147.6-51147.49" *)
  wire un1_main_basesoc_uart_tx_fifo_produce_ac0_0_TMR_1;
  (* src = "lattice_riscv.v:51147.6-51147.49" *)
  wire un1_main_basesoc_uart_tx_fifo_produce_ac0_0_TMR_2;
  (* src = "lattice_riscv.v:51084.6-51084.50" *)
  wire un1_main_basesoc_uart_tx_fifo_produce_axbxc0_TMR_0;
  (* src = "lattice_riscv.v:51084.6-51084.50" *)
  wire un1_main_basesoc_uart_tx_fifo_produce_axbxc0_TMR_1;
  (* src = "lattice_riscv.v:51084.6-51084.50" *)
  wire un1_main_basesoc_uart_tx_fifo_produce_axbxc0_TMR_2;
  (* src = "lattice_riscv.v:51085.6-51085.50" *)
  wire un1_main_basesoc_uart_tx_fifo_produce_axbxc1_TMR_0;
  (* src = "lattice_riscv.v:51085.6-51085.50" *)
  wire un1_main_basesoc_uart_tx_fifo_produce_axbxc1_TMR_1;
  (* src = "lattice_riscv.v:51085.6-51085.50" *)
  wire un1_main_basesoc_uart_tx_fifo_produce_axbxc1_TMR_2;
  (* src = "lattice_riscv.v:51086.6-51086.50" *)
  wire un1_main_basesoc_uart_tx_fifo_produce_axbxc2_TMR_0;
  (* src = "lattice_riscv.v:51086.6-51086.50" *)
  wire un1_main_basesoc_uart_tx_fifo_produce_axbxc2_TMR_1;
  (* src = "lattice_riscv.v:51086.6-51086.50" *)
  wire un1_main_basesoc_uart_tx_fifo_produce_axbxc2_TMR_2;
  (* src = "lattice_riscv.v:51089.6-51089.59" *)
  wire un1_main_basesoc_uart_tx_fifo_produce_axbxc3_N_13_mux_TMR_0;
  (* src = "lattice_riscv.v:51089.6-51089.59" *)
  wire un1_main_basesoc_uart_tx_fifo_produce_axbxc3_N_13_mux_TMR_1;
  (* src = "lattice_riscv.v:51089.6-51089.59" *)
  wire un1_main_basesoc_uart_tx_fifo_produce_axbxc3_N_13_mux_TMR_2;
  (* src = "lattice_riscv.v:51145.6-51145.57" *)
  wire un1_main_basesoc_uart_tx_fifo_produce_axbxc3_m6_e_0_TMR_0;
  (* src = "lattice_riscv.v:51145.6-51145.57" *)
  wire un1_main_basesoc_uart_tx_fifo_produce_axbxc3_m6_e_0_TMR_1;
  (* src = "lattice_riscv.v:51145.6-51145.57" *)
  wire un1_main_basesoc_uart_tx_fifo_produce_axbxc3_m6_e_0_TMR_2;
  (* src = "lattice_riscv.v:51146.6-51146.57" *)
  wire un1_main_basesoc_uart_tx_fifo_produce_axbxc3_m6_e_2_TMR_0;
  (* src = "lattice_riscv.v:51146.6-51146.57" *)
  wire un1_main_basesoc_uart_tx_fifo_produce_axbxc3_m6_e_2_TMR_1;
  (* src = "lattice_riscv.v:51146.6-51146.57" *)
  wire un1_main_basesoc_uart_tx_fifo_produce_axbxc3_m6_e_2_TMR_2;
  (* src = "lattice_riscv.v:51091.6-51091.57" *)
  wire un1_main_basesoc_uart_tx_fifo_produce_axbxc3_m6_e_3_TMR_0;
  (* src = "lattice_riscv.v:51091.6-51091.57" *)
  wire un1_main_basesoc_uart_tx_fifo_produce_axbxc3_m6_e_3_TMR_1;
  (* src = "lattice_riscv.v:51091.6-51091.57" *)
  wire un1_main_basesoc_uart_tx_fifo_produce_axbxc3_m6_e_3_TMR_2;
  (* src = "lattice_riscv.v:51164.6-51164.39" *)
  wire un1_main_crg_por_count_cry_0_0_S0_TMR_0;
  (* src = "lattice_riscv.v:51164.6-51164.39" *)
  wire un1_main_crg_por_count_cry_0_0_S0_TMR_1;
  (* src = "lattice_riscv.v:51164.6-51164.39" *)
  wire un1_main_crg_por_count_cry_0_0_S0_TMR_2;
  (* src = "lattice_riscv.v:51152.6-51152.39" *)
  wire un1_main_crg_por_count_cry_0_0_S1_TMR_0;
  (* src = "lattice_riscv.v:51152.6-51152.39" *)
  wire un1_main_crg_por_count_cry_0_0_S1_TMR_1;
  (* src = "lattice_riscv.v:51152.6-51152.39" *)
  wire un1_main_crg_por_count_cry_0_0_S1_TMR_2;
  (* src = "lattice_riscv.v:51011.6-51011.34" *)
  wire un1_main_crg_por_count_cry_0_TMR_0;
  (* src = "lattice_riscv.v:51011.6-51011.34" *)
  wire un1_main_crg_por_count_cry_0_TMR_1;
  (* src = "lattice_riscv.v:51011.6-51011.34" *)
  wire un1_main_crg_por_count_cry_0_TMR_2;
  (* src = "lattice_riscv.v:51016.6-51016.35" *)
  wire un1_main_crg_por_count_cry_10_TMR_0;
  (* src = "lattice_riscv.v:51016.6-51016.35" *)
  wire un1_main_crg_por_count_cry_10_TMR_1;
  (* src = "lattice_riscv.v:51016.6-51016.35" *)
  wire un1_main_crg_por_count_cry_10_TMR_2;
  (* src = "lattice_riscv.v:50854.6-50854.40" *)
  wire un1_main_crg_por_count_cry_11_0_S0_TMR_0;
  (* src = "lattice_riscv.v:50854.6-50854.40" *)
  wire un1_main_crg_por_count_cry_11_0_S0_TMR_1;
  (* src = "lattice_riscv.v:50854.6-50854.40" *)
  wire un1_main_crg_por_count_cry_11_0_S0_TMR_2;
  (* src = "lattice_riscv.v:50855.6-50855.40" *)
  wire un1_main_crg_por_count_cry_11_0_S1_TMR_0;
  (* src = "lattice_riscv.v:50855.6-50855.40" *)
  wire un1_main_crg_por_count_cry_11_0_S1_TMR_1;
  (* src = "lattice_riscv.v:50855.6-50855.40" *)
  wire un1_main_crg_por_count_cry_11_0_S1_TMR_2;
  (* src = "lattice_riscv.v:51017.6-51017.35" *)
  wire un1_main_crg_por_count_cry_12_TMR_0;
  (* src = "lattice_riscv.v:51017.6-51017.35" *)
  wire un1_main_crg_por_count_cry_12_TMR_1;
  (* src = "lattice_riscv.v:51017.6-51017.35" *)
  wire un1_main_crg_por_count_cry_12_TMR_2;
  (* src = "lattice_riscv.v:50856.6-50856.40" *)
  wire un1_main_crg_por_count_cry_13_0_S0_TMR_0;
  (* src = "lattice_riscv.v:50856.6-50856.40" *)
  wire un1_main_crg_por_count_cry_13_0_S0_TMR_1;
  (* src = "lattice_riscv.v:50856.6-50856.40" *)
  wire un1_main_crg_por_count_cry_13_0_S0_TMR_2;
  (* src = "lattice_riscv.v:50857.6-50857.40" *)
  wire un1_main_crg_por_count_cry_13_0_S1_TMR_0;
  (* src = "lattice_riscv.v:50857.6-50857.40" *)
  wire un1_main_crg_por_count_cry_13_0_S1_TMR_1;
  (* src = "lattice_riscv.v:50857.6-50857.40" *)
  wire un1_main_crg_por_count_cry_13_0_S1_TMR_2;
  (* src = "lattice_riscv.v:51018.6-51018.35" *)
  wire un1_main_crg_por_count_cry_14_TMR_0;
  (* src = "lattice_riscv.v:51018.6-51018.35" *)
  wire un1_main_crg_por_count_cry_14_TMR_1;
  (* src = "lattice_riscv.v:51018.6-51018.35" *)
  wire un1_main_crg_por_count_cry_14_TMR_2;
  (* src = "lattice_riscv.v:50844.6-50844.39" *)
  wire un1_main_crg_por_count_cry_1_0_S0_TMR_0;
  (* src = "lattice_riscv.v:50844.6-50844.39" *)
  wire un1_main_crg_por_count_cry_1_0_S0_TMR_1;
  (* src = "lattice_riscv.v:50844.6-50844.39" *)
  wire un1_main_crg_por_count_cry_1_0_S0_TMR_2;
  (* src = "lattice_riscv.v:50845.6-50845.39" *)
  wire un1_main_crg_por_count_cry_1_0_S1_TMR_0;
  (* src = "lattice_riscv.v:50845.6-50845.39" *)
  wire un1_main_crg_por_count_cry_1_0_S1_TMR_1;
  (* src = "lattice_riscv.v:50845.6-50845.39" *)
  wire un1_main_crg_por_count_cry_1_0_S1_TMR_2;
  (* src = "lattice_riscv.v:51012.6-51012.34" *)
  wire un1_main_crg_por_count_cry_2_TMR_0;
  (* src = "lattice_riscv.v:51012.6-51012.34" *)
  wire un1_main_crg_por_count_cry_2_TMR_1;
  (* src = "lattice_riscv.v:51012.6-51012.34" *)
  wire un1_main_crg_por_count_cry_2_TMR_2;
  (* src = "lattice_riscv.v:50846.6-50846.39" *)
  wire un1_main_crg_por_count_cry_3_0_S0_TMR_0;
  (* src = "lattice_riscv.v:50846.6-50846.39" *)
  wire un1_main_crg_por_count_cry_3_0_S0_TMR_1;
  (* src = "lattice_riscv.v:50846.6-50846.39" *)
  wire un1_main_crg_por_count_cry_3_0_S0_TMR_2;
  (* src = "lattice_riscv.v:50847.6-50847.39" *)
  wire un1_main_crg_por_count_cry_3_0_S1_TMR_0;
  (* src = "lattice_riscv.v:50847.6-50847.39" *)
  wire un1_main_crg_por_count_cry_3_0_S1_TMR_1;
  (* src = "lattice_riscv.v:50847.6-50847.39" *)
  wire un1_main_crg_por_count_cry_3_0_S1_TMR_2;
  (* src = "lattice_riscv.v:51013.6-51013.34" *)
  wire un1_main_crg_por_count_cry_4_TMR_0;
  (* src = "lattice_riscv.v:51013.6-51013.34" *)
  wire un1_main_crg_por_count_cry_4_TMR_1;
  (* src = "lattice_riscv.v:51013.6-51013.34" *)
  wire un1_main_crg_por_count_cry_4_TMR_2;
  (* src = "lattice_riscv.v:50848.6-50848.39" *)
  wire un1_main_crg_por_count_cry_5_0_S0_TMR_0;
  (* src = "lattice_riscv.v:50848.6-50848.39" *)
  wire un1_main_crg_por_count_cry_5_0_S0_TMR_1;
  (* src = "lattice_riscv.v:50848.6-50848.39" *)
  wire un1_main_crg_por_count_cry_5_0_S0_TMR_2;
  (* src = "lattice_riscv.v:50849.6-50849.39" *)
  wire un1_main_crg_por_count_cry_5_0_S1_TMR_0;
  (* src = "lattice_riscv.v:50849.6-50849.39" *)
  wire un1_main_crg_por_count_cry_5_0_S1_TMR_1;
  (* src = "lattice_riscv.v:50849.6-50849.39" *)
  wire un1_main_crg_por_count_cry_5_0_S1_TMR_2;
  (* src = "lattice_riscv.v:51014.6-51014.34" *)
  wire un1_main_crg_por_count_cry_6_TMR_0;
  (* src = "lattice_riscv.v:51014.6-51014.34" *)
  wire un1_main_crg_por_count_cry_6_TMR_1;
  (* src = "lattice_riscv.v:51014.6-51014.34" *)
  wire un1_main_crg_por_count_cry_6_TMR_2;
  (* src = "lattice_riscv.v:50850.6-50850.39" *)
  wire un1_main_crg_por_count_cry_7_0_S0_TMR_0;
  (* src = "lattice_riscv.v:50850.6-50850.39" *)
  wire un1_main_crg_por_count_cry_7_0_S0_TMR_1;
  (* src = "lattice_riscv.v:50850.6-50850.39" *)
  wire un1_main_crg_por_count_cry_7_0_S0_TMR_2;
  (* src = "lattice_riscv.v:50851.6-50851.39" *)
  wire un1_main_crg_por_count_cry_7_0_S1_TMR_0;
  (* src = "lattice_riscv.v:50851.6-50851.39" *)
  wire un1_main_crg_por_count_cry_7_0_S1_TMR_1;
  (* src = "lattice_riscv.v:50851.6-50851.39" *)
  wire un1_main_crg_por_count_cry_7_0_S1_TMR_2;
  (* src = "lattice_riscv.v:51015.6-51015.34" *)
  wire un1_main_crg_por_count_cry_8_TMR_0;
  (* src = "lattice_riscv.v:51015.6-51015.34" *)
  wire un1_main_crg_por_count_cry_8_TMR_1;
  (* src = "lattice_riscv.v:51015.6-51015.34" *)
  wire un1_main_crg_por_count_cry_8_TMR_2;
  (* src = "lattice_riscv.v:50852.6-50852.39" *)
  wire un1_main_crg_por_count_cry_9_0_S0_TMR_0;
  (* src = "lattice_riscv.v:50852.6-50852.39" *)
  wire un1_main_crg_por_count_cry_9_0_S0_TMR_1;
  (* src = "lattice_riscv.v:50852.6-50852.39" *)
  wire un1_main_crg_por_count_cry_9_0_S0_TMR_2;
  (* src = "lattice_riscv.v:50853.6-50853.39" *)
  wire un1_main_crg_por_count_cry_9_0_S1_TMR_0;
  (* src = "lattice_riscv.v:50853.6-50853.39" *)
  wire un1_main_crg_por_count_cry_9_0_S1_TMR_1;
  (* src = "lattice_riscv.v:50853.6-50853.39" *)
  wire un1_main_crg_por_count_cry_9_0_S1_TMR_2;
  (* src = "lattice_riscv.v:51166.6-51166.40" *)
  wire un1_main_crg_por_count_s_15_0_COUT_TMR_0;
  (* src = "lattice_riscv.v:51166.6-51166.40" *)
  wire un1_main_crg_por_count_s_15_0_COUT_TMR_1;
  (* src = "lattice_riscv.v:51166.6-51166.40" *)
  wire un1_main_crg_por_count_s_15_0_COUT_TMR_2;
  (* src = "lattice_riscv.v:50858.6-50858.38" *)
  wire un1_main_crg_por_count_s_15_0_S0_TMR_0;
  (* src = "lattice_riscv.v:50858.6-50858.38" *)
  wire un1_main_crg_por_count_s_15_0_S0_TMR_1;
  (* src = "lattice_riscv.v:50858.6-50858.38" *)
  wire un1_main_crg_por_count_s_15_0_S0_TMR_2;
  (* src = "lattice_riscv.v:51165.6-51165.38" *)
  wire un1_main_crg_por_count_s_15_0_S1_TMR_0;
  (* src = "lattice_riscv.v:51165.6-51165.38" *)
  wire un1_main_crg_por_count_s_15_0_S1_TMR_1;
  (* src = "lattice_riscv.v:51165.6-51165.38" *)
  wire un1_main_crg_por_count_s_15_0_S1_TMR_2;
  (* src = "lattice_riscv.v:50653.6-50653.29" *)
  wire un2_main_crg_por_done_1_TMR_0;
  (* src = "lattice_riscv.v:50653.6-50653.29" *)
  wire un2_main_crg_por_done_1_TMR_1;
  (* src = "lattice_riscv.v:50653.6-50653.29" *)
  wire un2_main_crg_por_done_1_TMR_2;
  (* src = "lattice_riscv.v:51092.6-51092.55" *)
  wire un3_main_basesoc_uart_tx_fifo_syncfifo_writable_i_TMR_0;
  (* src = "lattice_riscv.v:51092.6-51092.55" *)
  wire un3_main_basesoc_uart_tx_fifo_syncfifo_writable_i_TMR_1;
  (* src = "lattice_riscv.v:51092.6-51092.55" *)
  wire un3_main_basesoc_uart_tx_fifo_syncfifo_writable_i_TMR_2;
  (* src = "lattice_riscv.v:51162.6-51162.42" *)
  wire un5_main_basesoc_rx_phase_cry_0_0_S0_TMR_0;
  (* src = "lattice_riscv.v:51162.6-51162.42" *)
  wire un5_main_basesoc_rx_phase_cry_0_0_S0_TMR_1;
  (* src = "lattice_riscv.v:51162.6-51162.42" *)
  wire un5_main_basesoc_rx_phase_cry_0_0_S0_TMR_2;
  (* src = "lattice_riscv.v:51151.6-51151.42" *)
  wire un5_main_basesoc_rx_phase_cry_0_0_S1_TMR_0;
  (* src = "lattice_riscv.v:51151.6-51151.42" *)
  wire un5_main_basesoc_rx_phase_cry_0_0_S1_TMR_1;
  (* src = "lattice_riscv.v:51151.6-51151.42" *)
  wire un5_main_basesoc_rx_phase_cry_0_0_S1_TMR_2;
  (* src = "lattice_riscv.v:51019.6-51019.37" *)
  wire un5_main_basesoc_rx_phase_cry_0_TMR_0;
  (* src = "lattice_riscv.v:51019.6-51019.37" *)
  wire un5_main_basesoc_rx_phase_cry_0_TMR_1;
  (* src = "lattice_riscv.v:51019.6-51019.37" *)
  wire un5_main_basesoc_rx_phase_cry_0_TMR_2;
  (* src = "lattice_riscv.v:51024.6-51024.38" *)
  wire un5_main_basesoc_rx_phase_cry_10_TMR_0;
  (* src = "lattice_riscv.v:51024.6-51024.38" *)
  wire un5_main_basesoc_rx_phase_cry_10_TMR_1;
  (* src = "lattice_riscv.v:51024.6-51024.38" *)
  wire un5_main_basesoc_rx_phase_cry_10_TMR_2;
  (* src = "lattice_riscv.v:51025.6-51025.38" *)
  wire un5_main_basesoc_rx_phase_cry_12_TMR_0;
  (* src = "lattice_riscv.v:51025.6-51025.38" *)
  wire un5_main_basesoc_rx_phase_cry_12_TMR_1;
  (* src = "lattice_riscv.v:51025.6-51025.38" *)
  wire un5_main_basesoc_rx_phase_cry_12_TMR_2;
  (* src = "lattice_riscv.v:51026.6-51026.38" *)
  wire un5_main_basesoc_rx_phase_cry_14_TMR_0;
  (* src = "lattice_riscv.v:51026.6-51026.38" *)
  wire un5_main_basesoc_rx_phase_cry_14_TMR_1;
  (* src = "lattice_riscv.v:51026.6-51026.38" *)
  wire un5_main_basesoc_rx_phase_cry_14_TMR_2;
  (* src = "lattice_riscv.v:50827.6-50827.43" *)
  wire un5_main_basesoc_rx_phase_cry_15_0_S1_TMR_0;
  (* src = "lattice_riscv.v:50827.6-50827.43" *)
  wire un5_main_basesoc_rx_phase_cry_15_0_S1_TMR_1;
  (* src = "lattice_riscv.v:50827.6-50827.43" *)
  wire un5_main_basesoc_rx_phase_cry_15_0_S1_TMR_2;
  (* src = "lattice_riscv.v:51027.6-51027.38" *)
  wire un5_main_basesoc_rx_phase_cry_16_TMR_0;
  (* src = "lattice_riscv.v:51027.6-51027.38" *)
  wire un5_main_basesoc_rx_phase_cry_16_TMR_1;
  (* src = "lattice_riscv.v:51027.6-51027.38" *)
  wire un5_main_basesoc_rx_phase_cry_16_TMR_2;
  (* src = "lattice_riscv.v:51028.6-51028.38" *)
  wire un5_main_basesoc_rx_phase_cry_18_TMR_0;
  (* src = "lattice_riscv.v:51028.6-51028.38" *)
  wire un5_main_basesoc_rx_phase_cry_18_TMR_1;
  (* src = "lattice_riscv.v:51028.6-51028.38" *)
  wire un5_main_basesoc_rx_phase_cry_18_TMR_2;
  (* src = "lattice_riscv.v:50830.6-50830.43" *)
  wire un5_main_basesoc_rx_phase_cry_19_0_S0_TMR_0;
  (* src = "lattice_riscv.v:50830.6-50830.43" *)
  wire un5_main_basesoc_rx_phase_cry_19_0_S0_TMR_1;
  (* src = "lattice_riscv.v:50830.6-50830.43" *)
  wire un5_main_basesoc_rx_phase_cry_19_0_S0_TMR_2;
  (* src = "lattice_riscv.v:50831.6-50831.43" *)
  wire un5_main_basesoc_rx_phase_cry_19_0_S1_TMR_0;
  (* src = "lattice_riscv.v:50831.6-50831.43" *)
  wire un5_main_basesoc_rx_phase_cry_19_0_S1_TMR_1;
  (* src = "lattice_riscv.v:50831.6-50831.43" *)
  wire un5_main_basesoc_rx_phase_cry_19_0_S1_TMR_2;
  (* src = "lattice_riscv.v:51029.6-51029.38" *)
  wire un5_main_basesoc_rx_phase_cry_20_TMR_0;
  (* src = "lattice_riscv.v:51029.6-51029.38" *)
  wire un5_main_basesoc_rx_phase_cry_20_TMR_1;
  (* src = "lattice_riscv.v:51029.6-51029.38" *)
  wire un5_main_basesoc_rx_phase_cry_20_TMR_2;
  (* src = "lattice_riscv.v:51030.6-51030.38" *)
  wire un5_main_basesoc_rx_phase_cry_22_TMR_0;
  (* src = "lattice_riscv.v:51030.6-51030.38" *)
  wire un5_main_basesoc_rx_phase_cry_22_TMR_1;
  (* src = "lattice_riscv.v:51030.6-51030.38" *)
  wire un5_main_basesoc_rx_phase_cry_22_TMR_2;
  (* src = "lattice_riscv.v:50835.6-50835.43" *)
  wire un5_main_basesoc_rx_phase_cry_23_0_S1_TMR_0;
  (* src = "lattice_riscv.v:50835.6-50835.43" *)
  wire un5_main_basesoc_rx_phase_cry_23_0_S1_TMR_1;
  (* src = "lattice_riscv.v:50835.6-50835.43" *)
  wire un5_main_basesoc_rx_phase_cry_23_0_S1_TMR_2;
  (* src = "lattice_riscv.v:51031.6-51031.38" *)
  wire un5_main_basesoc_rx_phase_cry_24_TMR_0;
  (* src = "lattice_riscv.v:51031.6-51031.38" *)
  wire un5_main_basesoc_rx_phase_cry_24_TMR_1;
  (* src = "lattice_riscv.v:51031.6-51031.38" *)
  wire un5_main_basesoc_rx_phase_cry_24_TMR_2;
  (* src = "lattice_riscv.v:51032.6-51032.38" *)
  wire un5_main_basesoc_rx_phase_cry_26_TMR_0;
  (* src = "lattice_riscv.v:51032.6-51032.38" *)
  wire un5_main_basesoc_rx_phase_cry_26_TMR_1;
  (* src = "lattice_riscv.v:51032.6-51032.38" *)
  wire un5_main_basesoc_rx_phase_cry_26_TMR_2;
  (* src = "lattice_riscv.v:51033.6-51033.38" *)
  wire un5_main_basesoc_rx_phase_cry_28_TMR_0;
  (* src = "lattice_riscv.v:51033.6-51033.38" *)
  wire un5_main_basesoc_rx_phase_cry_28_TMR_1;
  (* src = "lattice_riscv.v:51033.6-51033.38" *)
  wire un5_main_basesoc_rx_phase_cry_28_TMR_2;
  (* src = "lattice_riscv.v:50840.6-50840.43" *)
  wire un5_main_basesoc_rx_phase_cry_29_0_S0_TMR_0;
  (* src = "lattice_riscv.v:50840.6-50840.43" *)
  wire un5_main_basesoc_rx_phase_cry_29_0_S0_TMR_1;
  (* src = "lattice_riscv.v:50840.6-50840.43" *)
  wire un5_main_basesoc_rx_phase_cry_29_0_S0_TMR_2;
  (* src = "lattice_riscv.v:50841.6-50841.43" *)
  wire un5_main_basesoc_rx_phase_cry_29_0_S1_TMR_0;
  (* src = "lattice_riscv.v:50841.6-50841.43" *)
  wire un5_main_basesoc_rx_phase_cry_29_0_S1_TMR_1;
  (* src = "lattice_riscv.v:50841.6-50841.43" *)
  wire un5_main_basesoc_rx_phase_cry_29_0_S1_TMR_2;
  (* src = "lattice_riscv.v:51020.6-51020.37" *)
  wire un5_main_basesoc_rx_phase_cry_2_TMR_0;
  (* src = "lattice_riscv.v:51020.6-51020.37" *)
  wire un5_main_basesoc_rx_phase_cry_2_TMR_1;
  (* src = "lattice_riscv.v:51020.6-51020.37" *)
  wire un5_main_basesoc_rx_phase_cry_2_TMR_2;
  (* src = "lattice_riscv.v:51034.6-51034.38" *)
  wire un5_main_basesoc_rx_phase_cry_30_TMR_0;
  (* src = "lattice_riscv.v:51034.6-51034.38" *)
  wire un5_main_basesoc_rx_phase_cry_30_TMR_1;
  (* src = "lattice_riscv.v:51034.6-51034.38" *)
  wire un5_main_basesoc_rx_phase_cry_30_TMR_2;
  (* src = "lattice_riscv.v:51163.6-51163.45" *)
  wire un5_main_basesoc_rx_phase_cry_31_0_COUT_TMR_0;
  (* src = "lattice_riscv.v:51163.6-51163.45" *)
  wire un5_main_basesoc_rx_phase_cry_31_0_COUT_TMR_1;
  (* src = "lattice_riscv.v:51163.6-51163.45" *)
  wire un5_main_basesoc_rx_phase_cry_31_0_COUT_TMR_2;
  (* src = "lattice_riscv.v:50842.6-50842.43" *)
  wire un5_main_basesoc_rx_phase_cry_31_0_S0_TMR_0;
  (* src = "lattice_riscv.v:50842.6-50842.43" *)
  wire un5_main_basesoc_rx_phase_cry_31_0_S0_TMR_1;
  (* src = "lattice_riscv.v:50842.6-50842.43" *)
  wire un5_main_basesoc_rx_phase_cry_31_0_S0_TMR_2;
  (* src = "lattice_riscv.v:50843.6-50843.38" *)
  wire un5_main_basesoc_rx_phase_cry_31_TMR_0;
  (* src = "lattice_riscv.v:50843.6-50843.38" *)
  wire un5_main_basesoc_rx_phase_cry_31_TMR_1;
  (* src = "lattice_riscv.v:50843.6-50843.38" *)
  wire un5_main_basesoc_rx_phase_cry_31_TMR_2;
  (* src = "lattice_riscv.v:51021.6-51021.37" *)
  wire un5_main_basesoc_rx_phase_cry_4_TMR_0;
  (* src = "lattice_riscv.v:51021.6-51021.37" *)
  wire un5_main_basesoc_rx_phase_cry_4_TMR_1;
  (* src = "lattice_riscv.v:51021.6-51021.37" *)
  wire un5_main_basesoc_rx_phase_cry_4_TMR_2;
  (* src = "lattice_riscv.v:51022.6-51022.37" *)
  wire un5_main_basesoc_rx_phase_cry_6_TMR_0;
  (* src = "lattice_riscv.v:51022.6-51022.37" *)
  wire un5_main_basesoc_rx_phase_cry_6_TMR_1;
  (* src = "lattice_riscv.v:51022.6-51022.37" *)
  wire un5_main_basesoc_rx_phase_cry_6_TMR_2;
  (* src = "lattice_riscv.v:51023.6-51023.37" *)
  wire un5_main_basesoc_rx_phase_cry_8_TMR_0;
  (* src = "lattice_riscv.v:51023.6-51023.37" *)
  wire un5_main_basesoc_rx_phase_cry_8_TMR_1;
  (* src = "lattice_riscv.v:51023.6-51023.37" *)
  wire un5_main_basesoc_rx_phase_cry_8_TMR_2;
  (* src = "lattice_riscv.v:51160.6-51160.42" *)
  wire un5_main_basesoc_tx_phase_cry_0_0_S0_TMR_0;
  (* src = "lattice_riscv.v:51160.6-51160.42" *)
  wire un5_main_basesoc_tx_phase_cry_0_0_S0_TMR_1;
  (* src = "lattice_riscv.v:51160.6-51160.42" *)
  wire un5_main_basesoc_tx_phase_cry_0_0_S0_TMR_2;
  (* src = "lattice_riscv.v:51150.6-51150.42" *)
  wire un5_main_basesoc_tx_phase_cry_0_0_S1_TMR_0;
  (* src = "lattice_riscv.v:51150.6-51150.42" *)
  wire un5_main_basesoc_tx_phase_cry_0_0_S1_TMR_1;
  (* src = "lattice_riscv.v:51150.6-51150.42" *)
  wire un5_main_basesoc_tx_phase_cry_0_0_S1_TMR_2;
  (* src = "lattice_riscv.v:51035.6-51035.37" *)
  wire un5_main_basesoc_tx_phase_cry_0_TMR_0;
  (* src = "lattice_riscv.v:51035.6-51035.37" *)
  wire un5_main_basesoc_tx_phase_cry_0_TMR_1;
  (* src = "lattice_riscv.v:51035.6-51035.37" *)
  wire un5_main_basesoc_tx_phase_cry_0_TMR_2;
  (* src = "lattice_riscv.v:51040.6-51040.38" *)
  wire un5_main_basesoc_tx_phase_cry_10_TMR_0;
  (* src = "lattice_riscv.v:51040.6-51040.38" *)
  wire un5_main_basesoc_tx_phase_cry_10_TMR_1;
  (* src = "lattice_riscv.v:51040.6-51040.38" *)
  wire un5_main_basesoc_tx_phase_cry_10_TMR_2;
  (* src = "lattice_riscv.v:50790.6-50790.43" *)
  wire un5_main_basesoc_tx_phase_cry_11_0_S0_TMR_0;
  (* src = "lattice_riscv.v:50790.6-50790.43" *)
  wire un5_main_basesoc_tx_phase_cry_11_0_S0_TMR_1;
  (* src = "lattice_riscv.v:50790.6-50790.43" *)
  wire un5_main_basesoc_tx_phase_cry_11_0_S0_TMR_2;
  (* src = "lattice_riscv.v:50791.6-50791.43" *)
  wire un5_main_basesoc_tx_phase_cry_11_0_S1_TMR_0;
  (* src = "lattice_riscv.v:50791.6-50791.43" *)
  wire un5_main_basesoc_tx_phase_cry_11_0_S1_TMR_1;
  (* src = "lattice_riscv.v:50791.6-50791.43" *)
  wire un5_main_basesoc_tx_phase_cry_11_0_S1_TMR_2;
  (* src = "lattice_riscv.v:51041.6-51041.38" *)
  wire un5_main_basesoc_tx_phase_cry_12_TMR_0;
  (* src = "lattice_riscv.v:51041.6-51041.38" *)
  wire un5_main_basesoc_tx_phase_cry_12_TMR_1;
  (* src = "lattice_riscv.v:51041.6-51041.38" *)
  wire un5_main_basesoc_tx_phase_cry_12_TMR_2;
  (* src = "lattice_riscv.v:50792.6-50792.43" *)
  wire un5_main_basesoc_tx_phase_cry_13_0_S0_TMR_0;
  (* src = "lattice_riscv.v:50792.6-50792.43" *)
  wire un5_main_basesoc_tx_phase_cry_13_0_S0_TMR_1;
  (* src = "lattice_riscv.v:50792.6-50792.43" *)
  wire un5_main_basesoc_tx_phase_cry_13_0_S0_TMR_2;
  (* src = "lattice_riscv.v:50793.6-50793.43" *)
  wire un5_main_basesoc_tx_phase_cry_13_0_S1_TMR_0;
  (* src = "lattice_riscv.v:50793.6-50793.43" *)
  wire un5_main_basesoc_tx_phase_cry_13_0_S1_TMR_1;
  (* src = "lattice_riscv.v:50793.6-50793.43" *)
  wire un5_main_basesoc_tx_phase_cry_13_0_S1_TMR_2;
  (* src = "lattice_riscv.v:51042.6-51042.38" *)
  wire un5_main_basesoc_tx_phase_cry_14_TMR_0;
  (* src = "lattice_riscv.v:51042.6-51042.38" *)
  wire un5_main_basesoc_tx_phase_cry_14_TMR_1;
  (* src = "lattice_riscv.v:51042.6-51042.38" *)
  wire un5_main_basesoc_tx_phase_cry_14_TMR_2;
  (* src = "lattice_riscv.v:50794.6-50794.43" *)
  wire un5_main_basesoc_tx_phase_cry_15_0_S0_TMR_0;
  (* src = "lattice_riscv.v:50794.6-50794.43" *)
  wire un5_main_basesoc_tx_phase_cry_15_0_S0_TMR_1;
  (* src = "lattice_riscv.v:50794.6-50794.43" *)
  wire un5_main_basesoc_tx_phase_cry_15_0_S0_TMR_2;
  (* src = "lattice_riscv.v:50795.6-50795.43" *)
  wire un5_main_basesoc_tx_phase_cry_15_0_S1_TMR_0;
  (* src = "lattice_riscv.v:50795.6-50795.43" *)
  wire un5_main_basesoc_tx_phase_cry_15_0_S1_TMR_1;
  (* src = "lattice_riscv.v:50795.6-50795.43" *)
  wire un5_main_basesoc_tx_phase_cry_15_0_S1_TMR_2;
  (* src = "lattice_riscv.v:51043.6-51043.38" *)
  wire un5_main_basesoc_tx_phase_cry_16_TMR_0;
  (* src = "lattice_riscv.v:51043.6-51043.38" *)
  wire un5_main_basesoc_tx_phase_cry_16_TMR_1;
  (* src = "lattice_riscv.v:51043.6-51043.38" *)
  wire un5_main_basesoc_tx_phase_cry_16_TMR_2;
  (* src = "lattice_riscv.v:50796.6-50796.43" *)
  wire un5_main_basesoc_tx_phase_cry_17_0_S0_TMR_0;
  (* src = "lattice_riscv.v:50796.6-50796.43" *)
  wire un5_main_basesoc_tx_phase_cry_17_0_S0_TMR_1;
  (* src = "lattice_riscv.v:50796.6-50796.43" *)
  wire un5_main_basesoc_tx_phase_cry_17_0_S0_TMR_2;
  (* src = "lattice_riscv.v:50797.6-50797.43" *)
  wire un5_main_basesoc_tx_phase_cry_17_0_S1_TMR_0;
  (* src = "lattice_riscv.v:50797.6-50797.43" *)
  wire un5_main_basesoc_tx_phase_cry_17_0_S1_TMR_1;
  (* src = "lattice_riscv.v:50797.6-50797.43" *)
  wire un5_main_basesoc_tx_phase_cry_17_0_S1_TMR_2;
  (* src = "lattice_riscv.v:51044.6-51044.38" *)
  wire un5_main_basesoc_tx_phase_cry_18_TMR_0;
  (* src = "lattice_riscv.v:51044.6-51044.38" *)
  wire un5_main_basesoc_tx_phase_cry_18_TMR_1;
  (* src = "lattice_riscv.v:51044.6-51044.38" *)
  wire un5_main_basesoc_tx_phase_cry_18_TMR_2;
  (* src = "lattice_riscv.v:50798.6-50798.43" *)
  wire un5_main_basesoc_tx_phase_cry_19_0_S0_TMR_0;
  (* src = "lattice_riscv.v:50798.6-50798.43" *)
  wire un5_main_basesoc_tx_phase_cry_19_0_S0_TMR_1;
  (* src = "lattice_riscv.v:50798.6-50798.43" *)
  wire un5_main_basesoc_tx_phase_cry_19_0_S0_TMR_2;
  (* src = "lattice_riscv.v:50799.6-50799.43" *)
  wire un5_main_basesoc_tx_phase_cry_19_0_S1_TMR_0;
  (* src = "lattice_riscv.v:50799.6-50799.43" *)
  wire un5_main_basesoc_tx_phase_cry_19_0_S1_TMR_1;
  (* src = "lattice_riscv.v:50799.6-50799.43" *)
  wire un5_main_basesoc_tx_phase_cry_19_0_S1_TMR_2;
  (* src = "lattice_riscv.v:50780.6-50780.42" *)
  wire un5_main_basesoc_tx_phase_cry_1_0_S0_TMR_0;
  (* src = "lattice_riscv.v:50780.6-50780.42" *)
  wire un5_main_basesoc_tx_phase_cry_1_0_S0_TMR_1;
  (* src = "lattice_riscv.v:50780.6-50780.42" *)
  wire un5_main_basesoc_tx_phase_cry_1_0_S0_TMR_2;
  (* src = "lattice_riscv.v:50781.6-50781.42" *)
  wire un5_main_basesoc_tx_phase_cry_1_0_S1_TMR_0;
  (* src = "lattice_riscv.v:50781.6-50781.42" *)
  wire un5_main_basesoc_tx_phase_cry_1_0_S1_TMR_1;
  (* src = "lattice_riscv.v:50781.6-50781.42" *)
  wire un5_main_basesoc_tx_phase_cry_1_0_S1_TMR_2;
  (* src = "lattice_riscv.v:51045.6-51045.38" *)
  wire un5_main_basesoc_tx_phase_cry_20_TMR_0;
  (* src = "lattice_riscv.v:51045.6-51045.38" *)
  wire un5_main_basesoc_tx_phase_cry_20_TMR_1;
  (* src = "lattice_riscv.v:51045.6-51045.38" *)
  wire un5_main_basesoc_tx_phase_cry_20_TMR_2;
  (* src = "lattice_riscv.v:50800.6-50800.43" *)
  wire un5_main_basesoc_tx_phase_cry_21_0_S0_TMR_0;
  (* src = "lattice_riscv.v:50800.6-50800.43" *)
  wire un5_main_basesoc_tx_phase_cry_21_0_S0_TMR_1;
  (* src = "lattice_riscv.v:50800.6-50800.43" *)
  wire un5_main_basesoc_tx_phase_cry_21_0_S0_TMR_2;
  (* src = "lattice_riscv.v:50801.6-50801.43" *)
  wire un5_main_basesoc_tx_phase_cry_21_0_S1_TMR_0;
  (* src = "lattice_riscv.v:50801.6-50801.43" *)
  wire un5_main_basesoc_tx_phase_cry_21_0_S1_TMR_1;
  (* src = "lattice_riscv.v:50801.6-50801.43" *)
  wire un5_main_basesoc_tx_phase_cry_21_0_S1_TMR_2;
  (* src = "lattice_riscv.v:51046.6-51046.38" *)
  wire un5_main_basesoc_tx_phase_cry_22_TMR_0;
  (* src = "lattice_riscv.v:51046.6-51046.38" *)
  wire un5_main_basesoc_tx_phase_cry_22_TMR_1;
  (* src = "lattice_riscv.v:51046.6-51046.38" *)
  wire un5_main_basesoc_tx_phase_cry_22_TMR_2;
  (* src = "lattice_riscv.v:50802.6-50802.43" *)
  wire un5_main_basesoc_tx_phase_cry_23_0_S0_TMR_0;
  (* src = "lattice_riscv.v:50802.6-50802.43" *)
  wire un5_main_basesoc_tx_phase_cry_23_0_S0_TMR_1;
  (* src = "lattice_riscv.v:50802.6-50802.43" *)
  wire un5_main_basesoc_tx_phase_cry_23_0_S0_TMR_2;
  (* src = "lattice_riscv.v:50803.6-50803.43" *)
  wire un5_main_basesoc_tx_phase_cry_23_0_S1_TMR_0;
  (* src = "lattice_riscv.v:50803.6-50803.43" *)
  wire un5_main_basesoc_tx_phase_cry_23_0_S1_TMR_1;
  (* src = "lattice_riscv.v:50803.6-50803.43" *)
  wire un5_main_basesoc_tx_phase_cry_23_0_S1_TMR_2;
  (* src = "lattice_riscv.v:51047.6-51047.38" *)
  wire un5_main_basesoc_tx_phase_cry_24_TMR_0;
  (* src = "lattice_riscv.v:51047.6-51047.38" *)
  wire un5_main_basesoc_tx_phase_cry_24_TMR_1;
  (* src = "lattice_riscv.v:51047.6-51047.38" *)
  wire un5_main_basesoc_tx_phase_cry_24_TMR_2;
  (* src = "lattice_riscv.v:50804.6-50804.43" *)
  wire un5_main_basesoc_tx_phase_cry_25_0_S0_TMR_0;
  (* src = "lattice_riscv.v:50804.6-50804.43" *)
  wire un5_main_basesoc_tx_phase_cry_25_0_S0_TMR_1;
  (* src = "lattice_riscv.v:50804.6-50804.43" *)
  wire un5_main_basesoc_tx_phase_cry_25_0_S0_TMR_2;
  (* src = "lattice_riscv.v:50805.6-50805.43" *)
  wire un5_main_basesoc_tx_phase_cry_25_0_S1_TMR_0;
  (* src = "lattice_riscv.v:50805.6-50805.43" *)
  wire un5_main_basesoc_tx_phase_cry_25_0_S1_TMR_1;
  (* src = "lattice_riscv.v:50805.6-50805.43" *)
  wire un5_main_basesoc_tx_phase_cry_25_0_S1_TMR_2;
  (* src = "lattice_riscv.v:51048.6-51048.38" *)
  wire un5_main_basesoc_tx_phase_cry_26_TMR_0;
  (* src = "lattice_riscv.v:51048.6-51048.38" *)
  wire un5_main_basesoc_tx_phase_cry_26_TMR_1;
  (* src = "lattice_riscv.v:51048.6-51048.38" *)
  wire un5_main_basesoc_tx_phase_cry_26_TMR_2;
  (* src = "lattice_riscv.v:50806.6-50806.43" *)
  wire un5_main_basesoc_tx_phase_cry_27_0_S0_TMR_0;
  (* src = "lattice_riscv.v:50806.6-50806.43" *)
  wire un5_main_basesoc_tx_phase_cry_27_0_S0_TMR_1;
  (* src = "lattice_riscv.v:50806.6-50806.43" *)
  wire un5_main_basesoc_tx_phase_cry_27_0_S0_TMR_2;
  (* src = "lattice_riscv.v:50807.6-50807.43" *)
  wire un5_main_basesoc_tx_phase_cry_27_0_S1_TMR_0;
  (* src = "lattice_riscv.v:50807.6-50807.43" *)
  wire un5_main_basesoc_tx_phase_cry_27_0_S1_TMR_1;
  (* src = "lattice_riscv.v:50807.6-50807.43" *)
  wire un5_main_basesoc_tx_phase_cry_27_0_S1_TMR_2;
  (* src = "lattice_riscv.v:51049.6-51049.38" *)
  wire un5_main_basesoc_tx_phase_cry_28_TMR_0;
  (* src = "lattice_riscv.v:51049.6-51049.38" *)
  wire un5_main_basesoc_tx_phase_cry_28_TMR_1;
  (* src = "lattice_riscv.v:51049.6-51049.38" *)
  wire un5_main_basesoc_tx_phase_cry_28_TMR_2;
  (* src = "lattice_riscv.v:50808.6-50808.43" *)
  wire un5_main_basesoc_tx_phase_cry_29_0_S0_TMR_0;
  (* src = "lattice_riscv.v:50808.6-50808.43" *)
  wire un5_main_basesoc_tx_phase_cry_29_0_S0_TMR_1;
  (* src = "lattice_riscv.v:50808.6-50808.43" *)
  wire un5_main_basesoc_tx_phase_cry_29_0_S0_TMR_2;
  (* src = "lattice_riscv.v:50809.6-50809.43" *)
  wire un5_main_basesoc_tx_phase_cry_29_0_S1_TMR_0;
  (* src = "lattice_riscv.v:50809.6-50809.43" *)
  wire un5_main_basesoc_tx_phase_cry_29_0_S1_TMR_1;
  (* src = "lattice_riscv.v:50809.6-50809.43" *)
  wire un5_main_basesoc_tx_phase_cry_29_0_S1_TMR_2;
  (* src = "lattice_riscv.v:51036.6-51036.37" *)
  wire un5_main_basesoc_tx_phase_cry_2_TMR_0;
  (* src = "lattice_riscv.v:51036.6-51036.37" *)
  wire un5_main_basesoc_tx_phase_cry_2_TMR_1;
  (* src = "lattice_riscv.v:51036.6-51036.37" *)
  wire un5_main_basesoc_tx_phase_cry_2_TMR_2;
  (* src = "lattice_riscv.v:51050.6-51050.38" *)
  wire un5_main_basesoc_tx_phase_cry_30_TMR_0;
  (* src = "lattice_riscv.v:51050.6-51050.38" *)
  wire un5_main_basesoc_tx_phase_cry_30_TMR_1;
  (* src = "lattice_riscv.v:51050.6-51050.38" *)
  wire un5_main_basesoc_tx_phase_cry_30_TMR_2;
  (* src = "lattice_riscv.v:51161.6-51161.45" *)
  wire un5_main_basesoc_tx_phase_cry_31_0_COUT_TMR_0;
  (* src = "lattice_riscv.v:51161.6-51161.45" *)
  wire un5_main_basesoc_tx_phase_cry_31_0_COUT_TMR_1;
  (* src = "lattice_riscv.v:51161.6-51161.45" *)
  wire un5_main_basesoc_tx_phase_cry_31_0_COUT_TMR_2;
  (* src = "lattice_riscv.v:50810.6-50810.43" *)
  wire un5_main_basesoc_tx_phase_cry_31_0_S0_TMR_0;
  (* src = "lattice_riscv.v:50810.6-50810.43" *)
  wire un5_main_basesoc_tx_phase_cry_31_0_S0_TMR_1;
  (* src = "lattice_riscv.v:50810.6-50810.43" *)
  wire un5_main_basesoc_tx_phase_cry_31_0_S0_TMR_2;
  (* src = "lattice_riscv.v:50811.6-50811.38" *)
  wire un5_main_basesoc_tx_phase_cry_31_TMR_0;
  (* src = "lattice_riscv.v:50811.6-50811.38" *)
  wire un5_main_basesoc_tx_phase_cry_31_TMR_1;
  (* src = "lattice_riscv.v:50811.6-50811.38" *)
  wire un5_main_basesoc_tx_phase_cry_31_TMR_2;
  (* src = "lattice_riscv.v:50782.6-50782.42" *)
  wire un5_main_basesoc_tx_phase_cry_3_0_S0_TMR_0;
  (* src = "lattice_riscv.v:50782.6-50782.42" *)
  wire un5_main_basesoc_tx_phase_cry_3_0_S0_TMR_1;
  (* src = "lattice_riscv.v:50782.6-50782.42" *)
  wire un5_main_basesoc_tx_phase_cry_3_0_S0_TMR_2;
  (* src = "lattice_riscv.v:50783.6-50783.42" *)
  wire un5_main_basesoc_tx_phase_cry_3_0_S1_TMR_0;
  (* src = "lattice_riscv.v:50783.6-50783.42" *)
  wire un5_main_basesoc_tx_phase_cry_3_0_S1_TMR_1;
  (* src = "lattice_riscv.v:50783.6-50783.42" *)
  wire un5_main_basesoc_tx_phase_cry_3_0_S1_TMR_2;
  (* src = "lattice_riscv.v:51037.6-51037.37" *)
  wire un5_main_basesoc_tx_phase_cry_4_TMR_0;
  (* src = "lattice_riscv.v:51037.6-51037.37" *)
  wire un5_main_basesoc_tx_phase_cry_4_TMR_1;
  (* src = "lattice_riscv.v:51037.6-51037.37" *)
  wire un5_main_basesoc_tx_phase_cry_4_TMR_2;
  (* src = "lattice_riscv.v:50784.6-50784.42" *)
  wire un5_main_basesoc_tx_phase_cry_5_0_S0_TMR_0;
  (* src = "lattice_riscv.v:50784.6-50784.42" *)
  wire un5_main_basesoc_tx_phase_cry_5_0_S0_TMR_1;
  (* src = "lattice_riscv.v:50784.6-50784.42" *)
  wire un5_main_basesoc_tx_phase_cry_5_0_S0_TMR_2;
  (* src = "lattice_riscv.v:50785.6-50785.42" *)
  wire un5_main_basesoc_tx_phase_cry_5_0_S1_TMR_0;
  (* src = "lattice_riscv.v:50785.6-50785.42" *)
  wire un5_main_basesoc_tx_phase_cry_5_0_S1_TMR_1;
  (* src = "lattice_riscv.v:50785.6-50785.42" *)
  wire un5_main_basesoc_tx_phase_cry_5_0_S1_TMR_2;
  (* src = "lattice_riscv.v:51038.6-51038.37" *)
  wire un5_main_basesoc_tx_phase_cry_6_TMR_0;
  (* src = "lattice_riscv.v:51038.6-51038.37" *)
  wire un5_main_basesoc_tx_phase_cry_6_TMR_1;
  (* src = "lattice_riscv.v:51038.6-51038.37" *)
  wire un5_main_basesoc_tx_phase_cry_6_TMR_2;
  (* src = "lattice_riscv.v:50786.6-50786.42" *)
  wire un5_main_basesoc_tx_phase_cry_7_0_S0_TMR_0;
  (* src = "lattice_riscv.v:50786.6-50786.42" *)
  wire un5_main_basesoc_tx_phase_cry_7_0_S0_TMR_1;
  (* src = "lattice_riscv.v:50786.6-50786.42" *)
  wire un5_main_basesoc_tx_phase_cry_7_0_S0_TMR_2;
  (* src = "lattice_riscv.v:50787.6-50787.42" *)
  wire un5_main_basesoc_tx_phase_cry_7_0_S1_TMR_0;
  (* src = "lattice_riscv.v:50787.6-50787.42" *)
  wire un5_main_basesoc_tx_phase_cry_7_0_S1_TMR_1;
  (* src = "lattice_riscv.v:50787.6-50787.42" *)
  wire un5_main_basesoc_tx_phase_cry_7_0_S1_TMR_2;
  (* src = "lattice_riscv.v:51039.6-51039.37" *)
  wire un5_main_basesoc_tx_phase_cry_8_TMR_0;
  (* src = "lattice_riscv.v:51039.6-51039.37" *)
  wire un5_main_basesoc_tx_phase_cry_8_TMR_1;
  (* src = "lattice_riscv.v:51039.6-51039.37" *)
  wire un5_main_basesoc_tx_phase_cry_8_TMR_2;
  (* src = "lattice_riscv.v:50788.6-50788.42" *)
  wire un5_main_basesoc_tx_phase_cry_9_0_S0_TMR_0;
  (* src = "lattice_riscv.v:50788.6-50788.42" *)
  wire un5_main_basesoc_tx_phase_cry_9_0_S0_TMR_1;
  (* src = "lattice_riscv.v:50788.6-50788.42" *)
  wire un5_main_basesoc_tx_phase_cry_9_0_S0_TMR_2;
  (* src = "lattice_riscv.v:50789.6-50789.42" *)
  wire un5_main_basesoc_tx_phase_cry_9_0_S1_TMR_0;
  (* src = "lattice_riscv.v:50789.6-50789.42" *)
  wire un5_main_basesoc_tx_phase_cry_9_0_S1_TMR_1;
  (* src = "lattice_riscv.v:50789.6-50789.42" *)
  wire un5_main_basesoc_tx_phase_cry_9_0_S1_TMR_2;
  (* src = "lattice_riscv.v:50450.8-50450.17" *)
  output user_led0;
  wire user_led0;
  wire user_led0_c_0_RED_VOTER_wire;
  (* src = "lattice_riscv.v:51188.6-51188.17" *)
  wire user_led0_c_TMR_0;
  (* src = "lattice_riscv.v:51188.6-51188.17" *)
  wire user_led0_c_TMR_1;
  (* src = "lattice_riscv.v:51188.6-51188.17" *)
  wire user_led0_c_TMR_2;
  (* src = "lattice_riscv.v:50451.8-50451.17" *)
  output user_led1;
  wire user_led1;
  (* src = "lattice_riscv.v:50460.8-50460.18" *)
  output user_led10;
  wire user_led10;
  wire user_led10_c_0_RED_VOTER_wire;
  (* src = "lattice_riscv.v:51198.6-51198.18" *)
  wire user_led10_c_TMR_0;
  (* src = "lattice_riscv.v:51198.6-51198.18" *)
  wire user_led10_c_TMR_1;
  (* src = "lattice_riscv.v:51198.6-51198.18" *)
  wire user_led10_c_TMR_2;
  (* src = "lattice_riscv.v:50461.8-50461.18" *)
  output user_led11;
  wire user_led11;
  wire user_led11_c_0_RED_VOTER_wire;
  (* src = "lattice_riscv.v:51199.6-51199.18" *)
  wire user_led11_c_TMR_0;
  (* src = "lattice_riscv.v:51199.6-51199.18" *)
  wire user_led11_c_TMR_1;
  (* src = "lattice_riscv.v:51199.6-51199.18" *)
  wire user_led11_c_TMR_2;
  (* src = "lattice_riscv.v:50462.8-50462.18" *)
  output user_led12;
  wire user_led12;
  wire user_led12_c_0_RED_VOTER_wire;
  (* src = "lattice_riscv.v:51200.6-51200.18" *)
  wire user_led12_c_TMR_0;
  (* src = "lattice_riscv.v:51200.6-51200.18" *)
  wire user_led12_c_TMR_1;
  (* src = "lattice_riscv.v:51200.6-51200.18" *)
  wire user_led12_c_TMR_2;
  (* src = "lattice_riscv.v:50463.8-50463.18" *)
  output user_led13;
  wire user_led13;
  wire user_led13_c_0_RED_VOTER_wire;
  (* src = "lattice_riscv.v:51201.6-51201.18" *)
  wire user_led13_c_TMR_0;
  (* src = "lattice_riscv.v:51201.6-51201.18" *)
  wire user_led13_c_TMR_1;
  (* src = "lattice_riscv.v:51201.6-51201.18" *)
  wire user_led13_c_TMR_2;
  wire user_led1_c_0_RED_VOTER_wire;
  (* src = "lattice_riscv.v:51189.6-51189.17" *)
  wire user_led1_c_TMR_0;
  (* src = "lattice_riscv.v:51189.6-51189.17" *)
  wire user_led1_c_TMR_1;
  (* src = "lattice_riscv.v:51189.6-51189.17" *)
  wire user_led1_c_TMR_2;
  (* src = "lattice_riscv.v:50452.8-50452.17" *)
  output user_led2;
  wire user_led2;
  wire user_led2_c_0_RED_VOTER_wire;
  (* src = "lattice_riscv.v:51190.6-51190.17" *)
  wire user_led2_c_TMR_0;
  (* src = "lattice_riscv.v:51190.6-51190.17" *)
  wire user_led2_c_TMR_1;
  (* src = "lattice_riscv.v:51190.6-51190.17" *)
  wire user_led2_c_TMR_2;
  (* src = "lattice_riscv.v:50453.8-50453.17" *)
  output user_led3;
  wire user_led3;
  wire user_led3_c_0_RED_VOTER_wire;
  (* src = "lattice_riscv.v:51191.6-51191.17" *)
  wire user_led3_c_TMR_0;
  (* src = "lattice_riscv.v:51191.6-51191.17" *)
  wire user_led3_c_TMR_1;
  (* src = "lattice_riscv.v:51191.6-51191.17" *)
  wire user_led3_c_TMR_2;
  (* src = "lattice_riscv.v:50454.8-50454.17" *)
  output user_led4;
  wire user_led4;
  wire user_led4_c_0_RED_VOTER_wire;
  (* src = "lattice_riscv.v:51192.6-51192.17" *)
  wire user_led4_c_TMR_0;
  (* src = "lattice_riscv.v:51192.6-51192.17" *)
  wire user_led4_c_TMR_1;
  (* src = "lattice_riscv.v:51192.6-51192.17" *)
  wire user_led4_c_TMR_2;
  (* src = "lattice_riscv.v:50455.8-50455.17" *)
  output user_led5;
  wire user_led5;
  wire user_led5_c_0_RED_VOTER_wire;
  (* src = "lattice_riscv.v:51193.6-51193.17" *)
  wire user_led5_c_TMR_0;
  (* src = "lattice_riscv.v:51193.6-51193.17" *)
  wire user_led5_c_TMR_1;
  (* src = "lattice_riscv.v:51193.6-51193.17" *)
  wire user_led5_c_TMR_2;
  (* src = "lattice_riscv.v:50456.8-50456.17" *)
  output user_led6;
  wire user_led6;
  wire user_led6_c_0_RED_VOTER_wire;
  (* src = "lattice_riscv.v:51194.6-51194.17" *)
  wire user_led6_c_TMR_0;
  (* src = "lattice_riscv.v:51194.6-51194.17" *)
  wire user_led6_c_TMR_1;
  (* src = "lattice_riscv.v:51194.6-51194.17" *)
  wire user_led6_c_TMR_2;
  (* src = "lattice_riscv.v:50457.8-50457.17" *)
  output user_led7;
  wire user_led7;
  wire user_led7_c_0_RED_VOTER_wire;
  (* src = "lattice_riscv.v:51195.6-51195.17" *)
  wire user_led7_c_TMR_0;
  (* src = "lattice_riscv.v:51195.6-51195.17" *)
  wire user_led7_c_TMR_1;
  (* src = "lattice_riscv.v:51195.6-51195.17" *)
  wire user_led7_c_TMR_2;
  (* src = "lattice_riscv.v:50458.8-50458.17" *)
  output user_led8;
  wire user_led8;
  wire user_led8_c_0_RED_VOTER_wire;
  (* src = "lattice_riscv.v:51196.6-51196.17" *)
  wire user_led8_c_TMR_0;
  (* src = "lattice_riscv.v:51196.6-51196.17" *)
  wire user_led8_c_TMR_1;
  (* src = "lattice_riscv.v:51196.6-51196.17" *)
  wire user_led8_c_TMR_2;
  (* src = "lattice_riscv.v:50459.8-50459.17" *)
  output user_led9;
  wire user_led9;
  wire user_led9_c_0_RED_VOTER_wire;
  (* src = "lattice_riscv.v:51197.6-51197.17" *)
  wire user_led9_c_TMR_0;
  (* src = "lattice_riscv.v:51197.6-51197.17" *)
  wire user_led9_c_TMR_1;
  (* src = "lattice_riscv.v:51197.6-51197.17" *)
  wire user_led9_c_TMR_2;
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:59319.11-59325.2" *)
  FD1P3BX FD1P3BX_1_TMR_0 (
    .CK(main_crg_clkout),
    .D(builder_rst10_TMR_0),
    .PD(gsrn_c_i_TMR_0),
    .Q(por_rst_TMR_0),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:59319.11-59325.2" *)
  FD1P3BX FD1P3BX_1_TMR_1 (
    .CK(main_crg_clkout),
    .D(builder_rst10_TMR_1),
    .PD(gsrn_c_i_TMR_1),
    .Q(por_rst_TMR_1),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:59319.11-59325.2" *)
  FD1P3BX FD1P3BX_1_TMR_2 (
    .CK(main_crg_clkout),
    .D(builder_rst10_TMR_2),
    .PD(gsrn_c_i_TMR_2),
    .Q(por_rst_TMR_2),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:59327.11-59333.2" *)
  FD1P3BX FD1P3BX_2_TMR_0 (
    .CK(sys_clk),
    .D(GND_0),
    .PD(un2_main_crg_por_done_1_TMR_0),
    .Q(builder_rst11_TMR_0),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:59327.11-59333.2" *)
  FD1P3BX FD1P3BX_2_TMR_1 (
    .CK(sys_clk),
    .D(GND_0),
    .PD(un2_main_crg_por_done_1_TMR_1),
    .Q(builder_rst11_TMR_1),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:59327.11-59333.2" *)
  FD1P3BX FD1P3BX_2_TMR_2 (
    .CK(sys_clk),
    .D(GND_0),
    .PD(un2_main_crg_por_done_1_TMR_2),
    .Q(builder_rst11_TMR_2),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:59335.11-59341.2" *)
  FD1P3BX FD1P3BX_3_TMR_0 (
    .CK(sys_clk),
    .D(builder_rst11_TMR_0),
    .PD(un2_main_crg_por_done_1_TMR_0),
    .Q(sys_rst_TMR_0),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:59335.11-59341.2" *)
  FD1P3BX FD1P3BX_3_TMR_1 (
    .CK(sys_clk),
    .D(builder_rst11_TMR_1),
    .PD(un2_main_crg_por_done_1_TMR_1),
    .Q(sys_rst_TMR_1),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:59335.11-59341.2" *)
  FD1P3BX FD1P3BX_3_TMR_2 (
    .CK(sys_clk),
    .D(builder_rst11_TMR_2),
    .PD(un2_main_crg_por_done_1_TMR_2),
    .Q(sys_rst_TMR_2),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:59311.11-59317.2" *)
  FD1P3BX FD1P3BX_TMR_0 (
    .CK(main_crg_clkout),
    .D(GND_0),
    .PD(gsrn_c_i_TMR_0),
    .Q(builder_rst10_TMR_0),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:59311.11-59317.2" *)
  FD1P3BX FD1P3BX_TMR_1 (
    .CK(main_crg_clkout),
    .D(GND_0),
    .PD(gsrn_c_i_TMR_1),
    .Q(builder_rst10_TMR_1),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:59311.11-59317.2" *)
  FD1P3BX FD1P3BX_TMR_2 (
    .CK(main_crg_clkout),
    .D(GND_0),
    .PD(gsrn_c_i_TMR_2),
    .Q(builder_rst10_TMR_2),
    .SP(VCC_TMR_2)
  );
  LUT4 GND_0_0_RED_VOTER (
    .A(GND_0),
    .B(GND_0),
    .C(GND_0),
    .D(1'h0),
    .Z(GND_0_0_RED_VOTER_wire)
  );
  defparam GND_0_0_RED_VOTER.INIT = "0xFCC0";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51259.7-51261.2" *)
  VLO GND_0_cZ_TMR_0 (
    .Z(GND_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51259.7-51261.2" *)
  VLO GND_0_cZ_TMR_1 (
    .Z(GND_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51259.7-51261.2" *)
  VLO GND_0_cZ_TMR_2 (
    .Z(GND_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51263.7-51266.2" *)
  GSR GSR_INST_TMR_0 (
    .CLK(NC0),
    .GSR_N(VCC_TMR_0)
  );
  defparam GSR_INST_TMR_0.SYNCMODE = "ASYNC";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51263.7-51266.2" *)
  GSR GSR_INST_TMR_1 (
    .CLK(NC0),
    .GSR_N(VCC_TMR_1)
  );
  defparam GSR_INST_TMR_1.SYNCMODE = "ASYNC";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51263.7-51266.2" *)
  GSR GSR_INST_TMR_2 (
    .CLK(NC0),
    .GSR_N(VCC_TMR_2)
  );
  defparam GSR_INST_TMR_2.SYNCMODE = "ASYNC";
  LUT4 N_103_0_RED_VOTER (
    .A(N_103_TMR_0),
    .B(N_103_TMR_1),
    .C(N_103_TMR_2),
    .D(1'h0),
    .Z(N_103_0_RED_VOTER_wire)
  );
  defparam N_103_0_RED_VOTER.INIT = "0xFCC0";
  LUT4 N_1209_i_0_RED_VOTER (
    .A(N_1209_i_TMR_0),
    .B(N_1209_i_TMR_1),
    .C(N_1209_i_TMR_2),
    .D(1'h0),
    .Z(N_1209_i_0_RED_VOTER_wire)
  );
  defparam N_1209_i_0_RED_VOTER.INIT = "0xFCC0";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:59429.8-59436.2" *)
  OSCA OSCA (
    .HFCLKCFG(HFCLKCFG),
    .HFCLKOUT(main_crg_clkout),
    .HFOUTEN(VCC_0_RED_VOTER_wire),
    .HFSDCOUT(HFSDCOUT),
    .HFSDSCEN(GND_0_0_RED_VOTER_wire),
    .LFCLKOUT(LFCLKOUT)
  );
  defparam OSCA.HF_CLK_DIV = "17";
  defparam OSCA.HF_OSC_EN = "ENABLED";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:59343.7-59399.2" *)
  PLL PLL_0 (
    .BINACT({ GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire }),
    .BINTEST({ GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire }),
    .CLKOP(sys_clk),
    .CLKOS(CLKOS),
    .CLKOS2(CLKOS2),
    .CLKOS3(CLKOS3),
    .CLKOS4(CLKOS4),
    .CLKOS5(builder_basesoc_clkfb),
    .CLKOUTDL(CLKOUTDL),
    .DIR(GND_0_0_RED_VOTER_wire),
    .DIRDEL(GND_0_0_RED_VOTER_wire),
    .DIRDELP1(GND_0_0_RED_VOTER_wire),
    .DIRSEL({ GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire }),
    .DYNROTATE(GND_0_0_RED_VOTER_wire),
    .ENCLKOP(GND_0_0_RED_VOTER_wire),
    .ENCLKOS(GND_0_0_RED_VOTER_wire),
    .ENCLKOS2(GND_0_0_RED_VOTER_wire),
    .ENCLKOS3(GND_0_0_RED_VOTER_wire),
    .ENCLKOS4(GND_0_0_RED_VOTER_wire),
    .ENCLKOS5(GND_0_0_RED_VOTER_wire),
    .FBKCK(builder_basesoc_clkfb),
    .GRAYACT({ GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire }),
    .GRAYTEST({ GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire }),
    .INTFBKOP(INTFBKOP),
    .INTFBKOS(INTFBKOS),
    .INTFBKOS2(INTFBKOS2),
    .INTFBKOS3(INTFBKOS3),
    .INTFBKOS4(INTFBKOS4),
    .INTFBKOS5(INTFBKOS5),
    .INTLOCK(INTLOCK),
    .LEGACY(GND_0_0_RED_VOTER_wire),
    .LEGRDYN(LEGRDYN),
    .LMMICLK(GND_0_0_RED_VOTER_wire),
    .LMMIOFFSET({ GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire }),
    .LMMIRDATA(LMMIRDATA),
    .LMMIRDATAVALID(LMMIRDATAVALID),
    .LMMIREADY(LMMIREADY),
    .LMMIREQUEST(GND_0_0_RED_VOTER_wire),
    .LMMIRESET_N(GND_0_0_RED_VOTER_wire),
    .LMMIWDATA({ GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire }),
    .LMMIWRRD_N(GND_0_0_RED_VOTER_wire),
    .LOADREG(GND_0_0_RED_VOTER_wire),
    .LOCK(main_crg_locked),
    .PFDDN(PFDDN),
    .PFDUP(PFDUP),
    .PLLPOWERDOWN_N(GND_0_0_RED_VOTER_wire),
    .PLLRESET(GND_0_0_RED_VOTER_wire),
    .REFCK(main_crg_clkout),
    .REFMUXCK(REFMUXCK),
    .REGQA(REGQA),
    .REGQB(REGQB),
    .REGQB1(REGQB1),
    .ROTDEL(GND_0_0_RED_VOTER_wire),
    .ROTDELP1(GND_0_0_RED_VOTER_wire),
    .STDBY(GND_0_0_RED_VOTER_wire)
  );
  defparam PLL_0.BW_CTL_BIAS = "0b1111";
  defparam PLL_0.CLKMUX_FB = "CMUX_CLKOS5";
  defparam PLL_0.CRIPPLE = "3P";
  defparam PLL_0.CSET = "8P";
  defparam PLL_0.DELA = "10";
  defparam PLL_0.DELF = "32";
  defparam PLL_0.DIVA = "10";
  defparam PLL_0.DIVF = "32";
  defparam PLL_0.ENCLK_CLKOP = "ENABLED";
  defparam PLL_0.ENCLK_CLKOS5 = "ENABLED";
  defparam PLL_0.FBK_INTEGER_MODE = "ENABLED";
  defparam PLL_0.FBK_MASK = "0b00000000";
  defparam PLL_0.FBK_MMD_DIG = "1";
  defparam PLL_0.IPI_CMP = "0b1100";
  defparam PLL_0.IPI_CMPN = "0b0011";
  defparam PLL_0.IPP_CTRL = "0b0110";
  defparam PLL_0.IPP_SEL = "0b1111";
  defparam PLL_0.KP_VCO = "0b00011";
  defparam PLL_0.PHIA = "0";
  defparam PLL_0.PLLPD_N = "USED";
  defparam PLL_0.PLLRESET_ENA = "ENABLED";
  defparam PLL_0.REF_INTEGER_MODE = "ENABLED";
  defparam PLL_0.REF_MMD_DIG = "1";
  defparam PLL_0.SEL_FBK = "FBKCLK5";
  defparam PLL_0.V2I_1V_EN = "ENABLED";
  defparam PLL_0.V2I_KVCO_SEL = "60";
  defparam PLL_0.V2I_PP_ICTRL = "0b11111";
  defparam PLL_0.V2I_PP_RES = "10K";
  (* ECC_BYTE_SEL = "BYTE_EN" *)
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:59279.38-59292.2" *)
  SP512K SP512K (
    .AD({ builder_array_muxed0_13_RED_VOTER_wire, builder_array_muxed0_12_RED_VOTER_wire, builder_array_muxed0_11_RED_VOTER_wire, builder_array_muxed0_10_RED_VOTER_wire, builder_array_muxed0_9_RED_VOTER_wire, builder_array_muxed0_8_RED_VOTER_wire, builder_array_muxed0_7_RED_VOTER_wire, builder_array_muxed0_6_RED_VOTER_wire, builder_array_muxed0_5_RED_VOTER_wire, builder_array_muxed0_4_RED_VOTER_wire, N_103_0_RED_VOTER_wire, builder_array_muxed0_2_RED_VOTER_wire, builder_array_muxed0_1_RED_VOTER_wire, builder_array_muxed0_0_RED_VOTER_wire }),
    .BYTEEN_N({ builder_array_muxed2_i_3_RED_VOTER_wire, builder_array_muxed2_i_2_RED_VOTER_wire, builder_array_muxed2_i_1_RED_VOTER_wire, builder_array_muxed2_i_0_RED_VOTER_wire }),
    .CE(VCC_0_RED_VOTER_wire),
    .CEOUT(GND_0_0_RED_VOTER_wire),
    .CLK(sys_clk),
    .CS(main_cs06_0_RED_VOTER_wire),
    .DI({ builder_array_muxed1_31_RED_VOTER_wire, builder_array_muxed1_30_RED_VOTER_wire, builder_array_muxed1_29_RED_VOTER_wire, builder_array_muxed1_28_RED_VOTER_wire, builder_array_muxed1_27_RED_VOTER_wire, builder_array_muxed1_26_RED_VOTER_wire, builder_array_muxed1_25_RED_VOTER_wire, builder_array_muxed1_24_RED_VOTER_wire, builder_array_muxed1_23_RED_VOTER_wire, builder_array_muxed1_22_RED_VOTER_wire, builder_array_muxed1_21_RED_VOTER_wire, builder_array_muxed1_20_RED_VOTER_wire, builder_array_muxed1_19_RED_VOTER_wire, builder_array_muxed1_18_RED_VOTER_wire, builder_array_muxed1_17_RED_VOTER_wire, builder_array_muxed1_16_RED_VOTER_wire, builder_array_muxed1_15_RED_VOTER_wire, builder_array_muxed1_14_RED_VOTER_wire, builder_array_muxed1_13_RED_VOTER_wire, builder_array_muxed1_12_RED_VOTER_wire, builder_array_muxed1_11_RED_VOTER_wire, builder_array_muxed1_10_RED_VOTER_wire, builder_array_muxed1_9_RED_VOTER_wire, builder_array_muxed1_8_RED_VOTER_wire, builder_array_muxed1_7_RED_VOTER_wire, builder_array_muxed1_6_RED_VOTER_wire, builder_array_muxed1_5_RED_VOTER_wire, builder_array_muxed1_4_RED_VOTER_wire, builder_array_muxed1_3_RED_VOTER_wire, builder_array_muxed1_2_RED_VOTER_wire, builder_array_muxed1_1_RED_VOTER_wire, builder_array_muxed1_0_RED_VOTER_wire }),
    .DO(main_dataout0),
    .ERRDECA(SP512K_ERRDECA),
    .ERRDECB(SP512K_ERRDECB),
    .RSTOUT(GND_0_0_RED_VOTER_wire),
    .WE(main_wren0_0_RED_VOTER_wire)
  );
  defparam SP512K.ECC_BYTE_SEL = "BYTE_EN";
  (* ECC_BYTE_SEL = "BYTE_EN" *)
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:59295.38-59308.2" *)
  SP512K SP512K_1 (
    .AD({ builder_array_muxed0_13_RED_VOTER_wire, builder_array_muxed0_12_RED_VOTER_wire, builder_array_muxed0_11_RED_VOTER_wire, builder_array_muxed0_10_RED_VOTER_wire, builder_array_muxed0_9_RED_VOTER_wire, builder_array_muxed0_8_RED_VOTER_wire, builder_array_muxed0_7_RED_VOTER_wire, builder_array_muxed0_6_RED_VOTER_wire, builder_array_muxed0_5_RED_VOTER_wire, builder_array_muxed0_4_RED_VOTER_wire, N_103_0_RED_VOTER_wire, builder_array_muxed0_2_RED_VOTER_wire, builder_array_muxed0_1_RED_VOTER_wire, builder_array_muxed0_0_RED_VOTER_wire }),
    .BYTEEN_N({ builder_array_muxed2_i_3_RED_VOTER_wire, builder_array_muxed2_i_2_RED_VOTER_wire, builder_array_muxed2_i_1_RED_VOTER_wire, builder_array_muxed2_i_0_RED_VOTER_wire }),
    .CE(VCC_0_RED_VOTER_wire),
    .CEOUT(GND_0_0_RED_VOTER_wire),
    .CLK(sys_clk),
    .CS(N_1209_i_0_RED_VOTER_wire),
    .DI({ builder_array_muxed1_31_RED_VOTER_wire, builder_array_muxed1_30_RED_VOTER_wire, builder_array_muxed1_29_RED_VOTER_wire, builder_array_muxed1_28_RED_VOTER_wire, builder_array_muxed1_27_RED_VOTER_wire, builder_array_muxed1_26_RED_VOTER_wire, builder_array_muxed1_25_RED_VOTER_wire, builder_array_muxed1_24_RED_VOTER_wire, builder_array_muxed1_23_RED_VOTER_wire, builder_array_muxed1_22_RED_VOTER_wire, builder_array_muxed1_21_RED_VOTER_wire, builder_array_muxed1_20_RED_VOTER_wire, builder_array_muxed1_19_RED_VOTER_wire, builder_array_muxed1_18_RED_VOTER_wire, builder_array_muxed1_17_RED_VOTER_wire, builder_array_muxed1_16_RED_VOTER_wire, builder_array_muxed1_15_RED_VOTER_wire, builder_array_muxed1_14_RED_VOTER_wire, builder_array_muxed1_13_RED_VOTER_wire, builder_array_muxed1_12_RED_VOTER_wire, builder_array_muxed1_11_RED_VOTER_wire, builder_array_muxed1_10_RED_VOTER_wire, builder_array_muxed1_9_RED_VOTER_wire, builder_array_muxed1_8_RED_VOTER_wire, builder_array_muxed1_7_RED_VOTER_wire, builder_array_muxed1_6_RED_VOTER_wire, builder_array_muxed1_5_RED_VOTER_wire, builder_array_muxed1_4_RED_VOTER_wire, builder_array_muxed1_3_RED_VOTER_wire, builder_array_muxed1_2_RED_VOTER_wire, builder_array_muxed1_1_RED_VOTER_wire, builder_array_muxed1_0_RED_VOTER_wire }),
    .DO(main_dataout1),
    .ERRDECA(SP512K_1_ERRDECA),
    .ERRDECB(SP512K_1_ERRDECB),
    .RSTOUT(GND_0_0_RED_VOTER_wire),
    .WE(main_wren1_0_RED_VOTER_wire)
  );
  defparam SP512K_1.ECC_BYTE_SEL = "BYTE_EN";
  LUT4 VCC_0_RED_VOTER (
    .A(VCC_TMR_0),
    .B(VCC_TMR_1),
    .C(VCC_TMR_2),
    .D(1'h0),
    .Z(VCC_0_RED_VOTER_wire)
  );
  defparam VCC_0_RED_VOTER.INIT = "0xFCC0";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51256.7-51258.2" *)
  VHI VCC_cZ_TMR_0 (
    .Z(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51256.7-51258.2" *)
  VHI VCC_cZ_TMR_1 (
    .Z(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51256.7-51258.2" *)
  VHI VCC_cZ_TMR_2 (
    .Z(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:59440.12-59629.2" *)
  VexRiscv VexRiscv (
    .CO0_0_TMR_0(CO0_0_TMR_0),
    .CO0_0_TMR_1(CO0_0_TMR_1),
    .CO0_0_TMR_2(CO0_0_TMR_2),
    .CO0_TMR_0(CO0_TMR_0),
    .CO0_TMR_1(CO0_TMR_1),
    .CO0_TMR_2(CO0_TMR_2),
    .N_100_TMR_0(N_100_TMR_0),
    .N_100_TMR_1(N_100_TMR_1),
    .N_100_TMR_2(N_100_TMR_2),
    .N_103_TMR_0(N_103_TMR_0),
    .N_103_TMR_1(N_103_TMR_1),
    .N_103_TMR_2(N_103_TMR_2),
    .N_110_TMR_0(N_110_TMR_0),
    .N_110_TMR_1(N_110_TMR_1),
    .N_110_TMR_2(N_110_TMR_2),
    .N_1209_i_TMR_0(N_1209_i_TMR_0),
    .N_1209_i_TMR_1(N_1209_i_TMR_1),
    .N_1209_i_TMR_2(N_1209_i_TMR_2),
    .N_120_i_TMR_0(N_120_i_TMR_0),
    .N_120_i_TMR_1(N_120_i_TMR_1),
    .N_120_i_TMR_2(N_120_i_TMR_2),
    .N_1210_i_TMR_0(N_1210_i_TMR_0),
    .N_1210_i_TMR_1(N_1210_i_TMR_1),
    .N_1210_i_TMR_2(N_1210_i_TMR_2),
    .N_1210_i_fast_TMR_0(N_1210_i_fast_TMR_0),
    .N_1210_i_fast_TMR_1(N_1210_i_fast_TMR_1),
    .N_1210_i_fast_TMR_2(N_1210_i_fast_TMR_2),
    .N_1210_i_rep1_TMR_0(N_1210_i_rep1_TMR_0),
    .N_1210_i_rep1_TMR_1(N_1210_i_rep1_TMR_1),
    .N_1210_i_rep1_TMR_2(N_1210_i_rep1_TMR_2),
    .N_1210_i_rep2_TMR_0(N_1210_i_rep2_TMR_0),
    .N_1210_i_rep2_TMR_1(N_1210_i_rep2_TMR_1),
    .N_1210_i_rep2_TMR_2(N_1210_i_rep2_TMR_2),
    .N_1218_i_TMR_0(N_1218_i_TMR_0),
    .N_1218_i_TMR_1(N_1218_i_TMR_1),
    .N_1218_i_TMR_2(N_1218_i_TMR_2),
    .N_1219_i_TMR_0(N_1219_i_TMR_0),
    .N_1219_i_TMR_1(N_1219_i_TMR_1),
    .N_1219_i_TMR_2(N_1219_i_TMR_2),
    .N_121_i_TMR_0(N_121_i_TMR_0),
    .N_121_i_TMR_1(N_121_i_TMR_1),
    .N_121_i_TMR_2(N_121_i_TMR_2),
    .N_123_i_TMR_0(N_123_i_TMR_0),
    .N_123_i_TMR_1(N_123_i_TMR_1),
    .N_123_i_TMR_2(N_123_i_TMR_2),
    .N_124_i_TMR_0(N_124_i_TMR_0),
    .N_124_i_TMR_1(N_124_i_TMR_1),
    .N_124_i_TMR_2(N_124_i_TMR_2),
    .N_136_TMR_0(N_136_TMR_0),
    .N_136_TMR_1(N_136_TMR_1),
    .N_136_TMR_2(N_136_TMR_2),
    .N_137_i_TMR_0(N_137_i_TMR_0),
    .N_137_i_TMR_1(N_137_i_TMR_1),
    .N_137_i_TMR_2(N_137_i_TMR_2),
    .N_148_TMR_0(N_148_TMR_0),
    .N_148_TMR_1(N_148_TMR_1),
    .N_148_TMR_2(N_148_TMR_2),
    .N_152_i_TMR_0(N_152_i_TMR_0),
    .N_152_i_TMR_1(N_152_i_TMR_1),
    .N_152_i_TMR_2(N_152_i_TMR_2),
    .N_167_TMR_0(N_167_TMR_0),
    .N_167_TMR_1(N_167_TMR_1),
    .N_167_TMR_2(N_167_TMR_2),
    .N_175_TMR_0(N_175_TMR_0),
    .N_175_TMR_1(N_175_TMR_1),
    .N_175_TMR_2(N_175_TMR_2),
    .N_20_TMR_0(N_20_TMR_0),
    .N_20_TMR_1(N_20_TMR_1),
    .N_20_TMR_2(N_20_TMR_2),
    .N_443_0_TMR_0(N_443_TMR_0),
    .N_443_0_TMR_1(N_443_TMR_1),
    .N_443_0_TMR_2(N_443_TMR_2),
    .N_792_0_TMR_0(N_792_TMR_0),
    .N_792_0_TMR_1(N_792_TMR_1),
    .N_792_0_TMR_2(N_792_TMR_2),
    .N_92_TMR_0(N_92_TMR_0),
    .N_92_TMR_1(N_92_TMR_1),
    .N_92_TMR_2(N_92_TMR_2),
    .builder_array_muxed0_TMR_0({ builder_array_muxed0_TMR_0[13:4], N_22657_TMR_0, builder_array_muxed0_TMR_0[2:0] }),
    .builder_array_muxed0_TMR_1({ builder_array_muxed0_TMR_1[13:4], N_22657_TMR_1, builder_array_muxed0_TMR_1[2:0] }),
    .builder_array_muxed0_TMR_2({ builder_array_muxed0_TMR_2[13:4], N_22657_TMR_2, builder_array_muxed0_TMR_2[2:0] }),
    .builder_array_muxed1_TMR_0(builder_array_muxed1_TMR_0),
    .builder_array_muxed1_TMR_1(builder_array_muxed1_TMR_1),
    .builder_array_muxed1_TMR_2(builder_array_muxed1_TMR_2),
    .builder_array_muxed2_i_TMR_0(builder_array_muxed2_i_TMR_0),
    .builder_array_muxed2_i_TMR_1(builder_array_muxed2_i_TMR_1),
    .builder_array_muxed2_i_TMR_2(builder_array_muxed2_i_TMR_2),
    .builder_basesoc_adr_TMR_0(builder_basesoc_adr_TMR_0),
    .builder_basesoc_adr_TMR_1(builder_basesoc_adr_TMR_1),
    .builder_basesoc_adr_TMR_2(builder_basesoc_adr_TMR_2),
    .builder_basesoc_next_state_1_sqmuxa_1_TMR_0(builder_basesoc_next_state_1_sqmuxa_1_TMR_0),
    .builder_basesoc_next_state_1_sqmuxa_1_TMR_1(builder_basesoc_next_state_1_sqmuxa_1_TMR_1),
    .builder_basesoc_next_state_1_sqmuxa_1_TMR_2(builder_basesoc_next_state_1_sqmuxa_1_TMR_2),
    .builder_basesoc_rs232phyrx_state_TMR_0(builder_basesoc_rs232phyrx_state_TMR_0),
    .builder_basesoc_rs232phyrx_state_TMR_1(builder_basesoc_rs232phyrx_state_TMR_1),
    .builder_basesoc_rs232phyrx_state_TMR_2(builder_basesoc_rs232phyrx_state_TMR_2),
    .builder_basesoc_rs232phytx_state_TMR_0(builder_basesoc_rs232phytx_state_TMR_0),
    .builder_basesoc_rs232phytx_state_TMR_1(builder_basesoc_rs232phytx_state_TMR_1),
    .builder_basesoc_rs232phytx_state_TMR_2(builder_basesoc_rs232phytx_state_TMR_2),
    .builder_basesoc_state_TMR_0(builder_basesoc_state_TMR_0),
    .builder_basesoc_state_TMR_1(builder_basesoc_state_TMR_1),
    .builder_basesoc_state_TMR_2(builder_basesoc_state_TMR_2),
    .builder_count_1_2_0_TMR_0(builder_count_1_2_TMR_0[6]),
    .builder_count_1_2_0_TMR_1(builder_count_1_2_TMR_1[6]),
    .builder_count_1_2_0_TMR_2(builder_count_1_2_TMR_2[6]),
    .builder_count_1_2_10_TMR_0(builder_count_1_2_TMR_0[16]),
    .builder_count_1_2_10_TMR_1(builder_count_1_2_TMR_1[16]),
    .builder_count_1_2_10_TMR_2(builder_count_1_2_TMR_2[16]),
    .builder_count_1_2_11_TMR_0(builder_count_1_2_TMR_0[17]),
    .builder_count_1_2_11_TMR_1(builder_count_1_2_TMR_1[17]),
    .builder_count_1_2_11_TMR_2(builder_count_1_2_TMR_2[17]),
    .builder_count_1_2_12_TMR_0(builder_count_1_2_TMR_0[18]),
    .builder_count_1_2_12_TMR_1(builder_count_1_2_TMR_1[18]),
    .builder_count_1_2_12_TMR_2(builder_count_1_2_TMR_2[18]),
    .builder_count_1_2_13_TMR_0(builder_count_1_2_TMR_0[19]),
    .builder_count_1_2_13_TMR_1(builder_count_1_2_TMR_1[19]),
    .builder_count_1_2_13_TMR_2(builder_count_1_2_TMR_2[19]),
    .builder_count_1_2_3_TMR_0(builder_count_1_2_TMR_0[9]),
    .builder_count_1_2_3_TMR_1(builder_count_1_2_TMR_1[9]),
    .builder_count_1_2_3_TMR_2(builder_count_1_2_TMR_2[9]),
    .builder_count_1_2_8_TMR_0(builder_count_1_2_TMR_0[14]),
    .builder_count_1_2_8_TMR_1(builder_count_1_2_TMR_1[14]),
    .builder_count_1_2_8_TMR_2(builder_count_1_2_TMR_2[14]),
    .builder_count_1_TMR_0(builder_count_1_TMR_0),
    .builder_count_1_TMR_1(builder_count_1_TMR_1),
    .builder_count_1_TMR_2(builder_count_1_TMR_2),
    .builder_count_1_cry_11_0_S1_TMR_0(builder_count_1_cry_11_0_S1_TMR_0),
    .builder_count_1_cry_11_0_S1_TMR_1(builder_count_1_cry_11_0_S1_TMR_1),
    .builder_count_1_cry_11_0_S1_TMR_2(builder_count_1_cry_11_0_S1_TMR_2),
    .builder_count_1_cry_15_0_S0_TMR_0(builder_count_1_cry_15_0_S0_TMR_0),
    .builder_count_1_cry_15_0_S0_TMR_1(builder_count_1_cry_15_0_S0_TMR_1),
    .builder_count_1_cry_15_0_S0_TMR_2(builder_count_1_cry_15_0_S0_TMR_2),
    .builder_count_r_0_TMR_0(builder_count_r_TMR_0[12]),
    .builder_count_r_0_TMR_1(builder_count_r_TMR_1[12]),
    .builder_count_r_0_TMR_2(builder_count_r_TMR_2[12]),
    .builder_count_r_3_TMR_0(builder_count_r_TMR_0[15]),
    .builder_count_r_3_TMR_1(builder_count_r_TMR_1[15]),
    .builder_count_r_3_TMR_2(builder_count_r_TMR_2[15]),
    .builder_csr_bankarray_csrbank0_reset0_re_1z_TMR_0(builder_csr_bankarray_csrbank0_reset0_re_TMR_0),
    .builder_csr_bankarray_csrbank0_reset0_re_1z_TMR_1(builder_csr_bankarray_csrbank0_reset0_re_TMR_1),
    .builder_csr_bankarray_csrbank0_reset0_re_1z_TMR_2(builder_csr_bankarray_csrbank0_reset0_re_TMR_2),
    .builder_csr_bankarray_csrbank0_scratch0_re_1z_TMR_0(builder_csr_bankarray_csrbank0_scratch0_re_TMR_0),
    .builder_csr_bankarray_csrbank0_scratch0_re_1z_TMR_1(builder_csr_bankarray_csrbank0_scratch0_re_TMR_1),
    .builder_csr_bankarray_csrbank0_scratch0_re_1z_TMR_2(builder_csr_bankarray_csrbank0_scratch0_re_TMR_2),
    .builder_csr_bankarray_csrbank1_out0_re_TMR_0(builder_csr_bankarray_csrbank1_out0_re_TMR_0),
    .builder_csr_bankarray_csrbank1_out0_re_TMR_1(builder_csr_bankarray_csrbank1_out0_re_TMR_1),
    .builder_csr_bankarray_csrbank1_out0_re_TMR_2(builder_csr_bankarray_csrbank1_out0_re_TMR_2),
    .builder_csr_bankarray_csrbank2_en0_re_1z_TMR_0(builder_csr_bankarray_csrbank2_en0_re_TMR_0),
    .builder_csr_bankarray_csrbank2_en0_re_1z_TMR_1(builder_csr_bankarray_csrbank2_en0_re_TMR_1),
    .builder_csr_bankarray_csrbank2_en0_re_1z_TMR_2(builder_csr_bankarray_csrbank2_en0_re_TMR_2),
    .builder_csr_bankarray_csrbank2_ev_enable0_re_1z_TMR_0(builder_csr_bankarray_csrbank2_ev_enable0_re_TMR_0),
    .builder_csr_bankarray_csrbank2_ev_enable0_re_1z_TMR_1(builder_csr_bankarray_csrbank2_ev_enable0_re_TMR_1),
    .builder_csr_bankarray_csrbank2_ev_enable0_re_1z_TMR_2(builder_csr_bankarray_csrbank2_ev_enable0_re_TMR_2),
    .builder_csr_bankarray_csrbank2_ev_pending_re_1z_TMR_0(builder_csr_bankarray_csrbank2_ev_pending_re_TMR_0),
    .builder_csr_bankarray_csrbank2_ev_pending_re_1z_TMR_1(builder_csr_bankarray_csrbank2_ev_pending_re_TMR_1),
    .builder_csr_bankarray_csrbank2_ev_pending_re_1z_TMR_2(builder_csr_bankarray_csrbank2_ev_pending_re_TMR_2),
    .builder_csr_bankarray_csrbank2_reload0_re_TMR_0(builder_csr_bankarray_csrbank2_reload0_re_TMR_0),
    .builder_csr_bankarray_csrbank2_reload0_re_TMR_1(builder_csr_bankarray_csrbank2_reload0_re_TMR_1),
    .builder_csr_bankarray_csrbank2_reload0_re_TMR_2(builder_csr_bankarray_csrbank2_reload0_re_TMR_2),
    .builder_csr_bankarray_csrbank2_update_value0_re_1z_TMR_0(builder_csr_bankarray_csrbank2_update_value0_re_TMR_0),
    .builder_csr_bankarray_csrbank2_update_value0_re_1z_TMR_1(builder_csr_bankarray_csrbank2_update_value0_re_TMR_1),
    .builder_csr_bankarray_csrbank2_update_value0_re_1z_TMR_2(builder_csr_bankarray_csrbank2_update_value0_re_TMR_2),
    .builder_csr_bankarray_csrbank3_ev_enable0_re_TMR_0(builder_csr_bankarray_csrbank3_ev_enable0_re_TMR_0),
    .builder_csr_bankarray_csrbank3_ev_enable0_re_TMR_1(builder_csr_bankarray_csrbank3_ev_enable0_re_TMR_1),
    .builder_csr_bankarray_csrbank3_ev_enable0_re_TMR_2(builder_csr_bankarray_csrbank3_ev_enable0_re_TMR_2),
    .builder_csr_bankarray_csrbank3_ev_pending_re_1z_TMR_0(builder_csr_bankarray_csrbank3_ev_pending_re_TMR_0),
    .builder_csr_bankarray_csrbank3_ev_pending_re_1z_TMR_1(builder_csr_bankarray_csrbank3_ev_pending_re_TMR_1),
    .builder_csr_bankarray_csrbank3_ev_pending_re_1z_TMR_2(builder_csr_bankarray_csrbank3_ev_pending_re_TMR_2),
    .builder_csr_bankarray_csrbank3_sel_TMR_0(builder_csr_bankarray_csrbank3_sel_TMR_0),
    .builder_csr_bankarray_csrbank3_sel_TMR_1(builder_csr_bankarray_csrbank3_sel_TMR_1),
    .builder_csr_bankarray_csrbank3_sel_TMR_2(builder_csr_bankarray_csrbank3_sel_TMR_2),
    .builder_csr_bankarray_dat_r_TMR_0({ builder_csr_bankarray_dat_r_TMR_0[7:6], N_22656, builder_csr_bankarray_dat_r_TMR_0[4:1] }),
    .builder_csr_bankarray_dat_r_TMR_1({ builder_csr_bankarray_dat_r_TMR_1[7:6], N_22656, builder_csr_bankarray_dat_r_TMR_1[4:1] }),
    .builder_csr_bankarray_dat_r_TMR_2({ builder_csr_bankarray_dat_r_TMR_2[7:6], N_22656, builder_csr_bankarray_dat_r_TMR_2[4:1] }),
    .builder_csr_bankarray_interface0_bank_bus_dat_r10_3_0_1z_TMR_0(\VexRiscv.builder_csr_bankarray_interface0_bank_bus_dat_r10_3_0_TMR_0 ),
    .builder_csr_bankarray_interface0_bank_bus_dat_r10_3_0_1z_TMR_1(\VexRiscv.builder_csr_bankarray_interface0_bank_bus_dat_r10_3_0_TMR_1 ),
    .builder_csr_bankarray_interface0_bank_bus_dat_r10_3_0_1z_TMR_2(\VexRiscv.builder_csr_bankarray_interface0_bank_bus_dat_r10_3_0_TMR_2 ),
    .builder_csr_bankarray_interface0_bank_bus_dat_r8_0_1z_TMR_0(\VexRiscv.builder_csr_bankarray_interface0_bank_bus_dat_r8_0_TMR_0 ),
    .builder_csr_bankarray_interface0_bank_bus_dat_r8_0_1z_TMR_1(\VexRiscv.builder_csr_bankarray_interface0_bank_bus_dat_r8_0_TMR_1 ),
    .builder_csr_bankarray_interface0_bank_bus_dat_r8_0_1z_TMR_2(\VexRiscv.builder_csr_bankarray_interface0_bank_bus_dat_r8_0_TMR_2 ),
    .builder_csr_bankarray_interface0_bank_bus_dat_r8_6_RNIG6FO8_TMR_0(builder_csr_bankarray_interface0_bank_bus_dat_r8_6_RNIG6FO8_TMR_0),
    .builder_csr_bankarray_interface0_bank_bus_dat_r8_6_RNIG6FO8_TMR_1(builder_csr_bankarray_interface0_bank_bus_dat_r8_6_RNIG6FO8_TMR_1),
    .builder_csr_bankarray_interface0_bank_bus_dat_r8_6_RNIG6FO8_TMR_2(builder_csr_bankarray_interface0_bank_bus_dat_r8_6_RNIG6FO8_TMR_2),
    .builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_0({ builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_0[31:2], N_22659_TMR_0, builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_0[0] }),
    .builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_1({ builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_1[31:2], N_22659_TMR_1, builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_1[0] }),
    .builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_2({ builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_2[31:2], N_22659_TMR_2, builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_2[0] }),
    .builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_0(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_0 ),
    .builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_1(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_1 ),
    .builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_2(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_2 ),
    .builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_0({ builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_0[31:2], N_22658, builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_0[0] }),
    .builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_1({ builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_1[31:2], N_22658, builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_1[0] }),
    .builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_2({ builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_2[31:2], N_22658, builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_2[0] }),
    .builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_0(builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_0),
    .builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_1(builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_1),
    .builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_2(builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_2),
    .builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_0(builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_0),
    .builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_1(builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_1),
    .builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_2(builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_2),
    .builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_0(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_0),
    .builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_1(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_1),
    .builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_2(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_2),
    .builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_0(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_0),
    .builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_1(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_1),
    .builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_2(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_2),
    .builder_csr_bankarray_interface3_bank_bus_dat_r_0_sqmuxa_1z_TMR_0(builder_csr_bankarray_interface3_bank_bus_dat_r_0_sqmuxa_TMR_0),
    .builder_csr_bankarray_interface3_bank_bus_dat_r_0_sqmuxa_1z_TMR_1(builder_csr_bankarray_interface3_bank_bus_dat_r_0_sqmuxa_TMR_1),
    .builder_csr_bankarray_interface3_bank_bus_dat_r_0_sqmuxa_1z_TMR_2(builder_csr_bankarray_interface3_bank_bus_dat_r_0_sqmuxa_TMR_2),
    .builder_csr_bankarray_interface3_bank_bus_dat_r_0_sqmuxa_i_TMR_0(builder_csr_bankarray_interface3_bank_bus_dat_r_0_sqmuxa_i_TMR_0),
    .builder_csr_bankarray_interface3_bank_bus_dat_r_0_sqmuxa_i_TMR_1(builder_csr_bankarray_interface3_bank_bus_dat_r_0_sqmuxa_i_TMR_1),
    .builder_csr_bankarray_interface3_bank_bus_dat_r_0_sqmuxa_i_TMR_2(builder_csr_bankarray_interface3_bank_bus_dat_r_0_sqmuxa_i_TMR_2),
    .builder_csr_bankarray_interface3_bank_bus_dat_r_11_TMR_0(builder_csr_bankarray_interface3_bank_bus_dat_r_11_TMR_0),
    .builder_csr_bankarray_interface3_bank_bus_dat_r_11_TMR_1(builder_csr_bankarray_interface3_bank_bus_dat_r_11_TMR_1),
    .builder_csr_bankarray_interface3_bank_bus_dat_r_11_TMR_2(builder_csr_bankarray_interface3_bank_bus_dat_r_11_TMR_2),
    .builder_csr_bankarray_interface3_bank_bus_dat_r_TMR_0(builder_csr_bankarray_interface3_bank_bus_dat_r_TMR_0),
    .builder_csr_bankarray_interface3_bank_bus_dat_r_TMR_1(builder_csr_bankarray_interface3_bank_bus_dat_r_TMR_1),
    .builder_csr_bankarray_interface3_bank_bus_dat_r_TMR_2(builder_csr_bankarray_interface3_bank_bus_dat_r_TMR_2),
    .builder_csr_bankarray_sel_r_TMR_0(builder_csr_bankarray_sel_r_TMR_0),
    .builder_csr_bankarray_sel_r_TMR_1(builder_csr_bankarray_sel_r_TMR_1),
    .builder_csr_bankarray_sel_r_TMR_2(builder_csr_bankarray_sel_r_TMR_2),
    .builder_csr_bankarray_sel_r_r_0_a2_TMR_0(builder_csr_bankarray_sel_r_r_0_a2_TMR_0),
    .builder_csr_bankarray_sel_r_r_0_a2_TMR_1(builder_csr_bankarray_sel_r_r_0_a2_TMR_1),
    .builder_csr_bankarray_sel_r_r_0_a2_TMR_2(builder_csr_bankarray_sel_r_r_0_a2_TMR_2),
    .builder_grant_TMR_0(builder_grant_TMR_0),
    .builder_grant_TMR_1(builder_grant_TMR_1),
    .builder_grant_TMR_2(builder_grant_TMR_2),
    .builder_grant_fast_TMR_0(builder_grant_fast_TMR_0),
    .builder_grant_fast_TMR_1(builder_grant_fast_TMR_1),
    .builder_grant_fast_TMR_2(builder_grant_fast_TMR_2),
    .builder_grant_rep1_TMR_0(builder_grant_rep1_TMR_0),
    .builder_grant_rep1_TMR_1(builder_grant_rep1_TMR_1),
    .builder_grant_rep1_TMR_2(builder_grant_rep1_TMR_2),
    .builder_grant_rep2_TMR_0(builder_grant_rep2_TMR_0),
    .builder_grant_rep2_TMR_1(builder_grant_rep2_TMR_1),
    .builder_grant_rep2_TMR_2(builder_grant_rep2_TMR_2),
    .builder_regs1_TMR_0(builder_regs1_TMR_0),
    .builder_regs1_TMR_1(builder_regs1_TMR_1),
    .builder_regs1_TMR_2(builder_regs1_TMR_2),
    .builder_slave_sel_2_0_TMR_0(builder_slave_sel_2_TMR_0),
    .builder_slave_sel_2_0_TMR_1(builder_slave_sel_2_TMR_1),
    .builder_slave_sel_2_0_TMR_2(builder_slave_sel_2_TMR_2),
    .builder_slave_sel_r_TMR_0(builder_slave_sel_r_TMR_0),
    .builder_slave_sel_r_TMR_1(builder_slave_sel_r_TMR_1),
    .builder_slave_sel_r_TMR_2(builder_slave_sel_r_TMR_2),
    .builder_slave_sel_r_r_0_a2_0_TMR_0(builder_slave_sel_r_r_0_a2_TMR_0),
    .builder_slave_sel_r_r_0_a2_0_TMR_1(builder_slave_sel_r_r_0_a2_TMR_1),
    .builder_slave_sel_r_r_0_a2_0_TMR_2(builder_slave_sel_r_r_0_a2_TMR_2),
    .builder_slave_sel_r_r_0_a2_0_out_TMR_0(\VexRiscv.IBusCachedPlugin_cache.builder_slave_sel_r_r_0_a2_0_out_TMR_0 ),
    .builder_slave_sel_r_r_0_a2_0_out_TMR_1(\VexRiscv.IBusCachedPlugin_cache.builder_slave_sel_r_r_0_a2_0_out_TMR_1 ),
    .builder_slave_sel_r_r_0_a2_0_out_TMR_2(\VexRiscv.IBusCachedPlugin_cache.builder_slave_sel_r_r_0_a2_0_out_TMR_2 ),
    .builder_wait_TMR_0(builder_wait_TMR_0),
    .builder_wait_TMR_1(builder_wait_TMR_1),
    .builder_wait_TMR_2(builder_wait_TMR_2),
    .dsp_join_kb_0_TMR_0(dsp_join_kb_0_TMR_0),
    .dsp_join_kb_0_TMR_1(dsp_join_kb_0_TMR_1),
    .dsp_join_kb_0_TMR_2(dsp_join_kb_0_TMR_2),
    .dsp_join_kb_25_TMR_0(dsp_join_kb_25_TMR_0),
    .dsp_join_kb_25_TMR_1(dsp_join_kb_25_TMR_1),
    .dsp_join_kb_25_TMR_2(dsp_join_kb_25_TMR_2),
    .dsp_join_kb_TMR_0(dsp_join_kb_TMR_0),
    .dsp_join_kb_TMR_1(dsp_join_kb_TMR_1),
    .dsp_join_kb_TMR_2(dsp_join_kb_TMR_2),
    .dsp_split_kb_0_TMR_0(dsp_split_kb_0_TMR_0),
    .dsp_split_kb_0_TMR_1(dsp_split_kb_0_TMR_1),
    .dsp_split_kb_0_TMR_2(dsp_split_kb_0_TMR_2),
    .dsp_split_kb_1_TMR_0(dsp_split_kb_1_TMR_0),
    .dsp_split_kb_1_TMR_1(dsp_split_kb_1_TMR_1),
    .dsp_split_kb_1_TMR_2(dsp_split_kb_1_TMR_2),
    .m71_TMR_0(m71_TMR_0),
    .m71_TMR_1(m71_TMR_1),
    .m71_TMR_2(m71_TMR_2),
    .main_basesoc_bus_errors_0_sqmuxa_TMR_0(main_basesoc_bus_errors_0_sqmuxa_TMR_0),
    .main_basesoc_bus_errors_0_sqmuxa_TMR_1(main_basesoc_bus_errors_0_sqmuxa_TMR_1),
    .main_basesoc_bus_errors_0_sqmuxa_TMR_2(main_basesoc_bus_errors_0_sqmuxa_TMR_2),
    .main_basesoc_ram_bus_ack_TMR_0(main_basesoc_ram_bus_ack_TMR_0),
    .main_basesoc_ram_bus_ack_TMR_1(main_basesoc_ram_bus_ack_TMR_1),
    .main_basesoc_ram_bus_ack_TMR_2(main_basesoc_ram_bus_ack_TMR_2),
    .main_basesoc_ram_bus_ack_r_TMR_0(main_basesoc_ram_bus_ack_r_TMR_0),
    .main_basesoc_ram_bus_ack_r_TMR_1(main_basesoc_ram_bus_ack_r_TMR_1),
    .main_basesoc_ram_bus_ack_r_TMR_2(main_basesoc_ram_bus_ack_r_TMR_2),
    .main_basesoc_reset_re_TMR_0(main_basesoc_reset_re_TMR_0),
    .main_basesoc_reset_re_TMR_1(main_basesoc_reset_re_TMR_1),
    .main_basesoc_reset_re_TMR_2(main_basesoc_reset_re_TMR_2),
    .main_basesoc_reset_storage_0_sqmuxa_1z_TMR_0(main_basesoc_reset_storage_0_sqmuxa_TMR_0),
    .main_basesoc_reset_storage_0_sqmuxa_1z_TMR_1(main_basesoc_reset_storage_0_sqmuxa_TMR_1),
    .main_basesoc_reset_storage_0_sqmuxa_1z_TMR_2(main_basesoc_reset_storage_0_sqmuxa_TMR_2),
    .main_basesoc_reset_storage_TMR_0(main_basesoc_reset_storage_TMR_0),
    .main_basesoc_reset_storage_TMR_1(main_basesoc_reset_storage_TMR_1),
    .main_basesoc_reset_storage_TMR_2(main_basesoc_reset_storage_TMR_2),
    .main_basesoc_rx_count_TMR_0(main_basesoc_rx_count_TMR_0),
    .main_basesoc_rx_count_TMR_1(main_basesoc_rx_count_TMR_1),
    .main_basesoc_rx_count_TMR_2(main_basesoc_rx_count_TMR_2),
    .main_basesoc_rx_count_rs232phyrx_next_value0_TMR_0(main_basesoc_rx_count_rs232phyrx_next_value0_TMR_0),
    .main_basesoc_rx_count_rs232phyrx_next_value0_TMR_1(main_basesoc_rx_count_rs232phyrx_next_value0_TMR_1),
    .main_basesoc_rx_count_rs232phyrx_next_value0_TMR_2(main_basesoc_rx_count_rs232phyrx_next_value0_TMR_2),
    .main_basesoc_rx_count_rs232phyrx_next_value_ce0_TMR_0(main_basesoc_rx_count_rs232phyrx_next_value_ce0_TMR_0),
    .main_basesoc_rx_count_rs232phyrx_next_value_ce0_TMR_1(main_basesoc_rx_count_rs232phyrx_next_value_ce0_TMR_1),
    .main_basesoc_rx_count_rs232phyrx_next_value_ce0_TMR_2(main_basesoc_rx_count_rs232phyrx_next_value_ce0_TMR_2),
    .main_basesoc_rx_data_TMR_0(main_basesoc_rx_data_TMR_0),
    .main_basesoc_rx_data_TMR_1(main_basesoc_rx_data_TMR_1),
    .main_basesoc_rx_data_TMR_2(main_basesoc_rx_data_TMR_2),
    .main_basesoc_rx_data_rs232phyrx_next_value1_0_sqmuxa_TMR_0(main_basesoc_rx_data_rs232phyrx_next_value1_0_sqmuxa_TMR_0),
    .main_basesoc_rx_data_rs232phyrx_next_value1_0_sqmuxa_TMR_1(main_basesoc_rx_data_rs232phyrx_next_value1_0_sqmuxa_TMR_1),
    .main_basesoc_rx_data_rs232phyrx_next_value1_0_sqmuxa_TMR_2(main_basesoc_rx_data_rs232phyrx_next_value1_0_sqmuxa_TMR_2),
    .main_basesoc_rx_rx_d_TMR_0(main_basesoc_rx_rx_d_TMR_0),
    .main_basesoc_rx_rx_d_TMR_1(main_basesoc_rx_rx_d_TMR_1),
    .main_basesoc_rx_rx_d_TMR_2(main_basesoc_rx_rx_d_TMR_2),
    .main_basesoc_rx_source_payload_data_TMR_0(main_basesoc_rx_source_payload_data_TMR_0),
    .main_basesoc_rx_source_payload_data_TMR_1(main_basesoc_rx_source_payload_data_TMR_1),
    .main_basesoc_rx_source_payload_data_TMR_2(main_basesoc_rx_source_payload_data_TMR_2),
    .main_basesoc_rx_tick_0_TMR_0(main_basesoc_rx_tick_0_TMR_0),
    .main_basesoc_rx_tick_0_TMR_1(main_basesoc_rx_tick_0_TMR_1),
    .main_basesoc_rx_tick_0_TMR_2(main_basesoc_rx_tick_0_TMR_2),
    .main_basesoc_rx_tick_TMR_0(main_basesoc_rx_tick_TMR_0),
    .main_basesoc_rx_tick_TMR_1(main_basesoc_rx_tick_TMR_1),
    .main_basesoc_rx_tick_TMR_2(main_basesoc_rx_tick_TMR_2),
    .main_basesoc_scratch_storage_TMR_0(main_basesoc_scratch_storage_TMR_0),
    .main_basesoc_scratch_storage_TMR_1(main_basesoc_scratch_storage_TMR_1),
    .main_basesoc_scratch_storage_TMR_2(main_basesoc_scratch_storage_TMR_2),
    .main_basesoc_serial_tx_rs232phytx_next_value1_1_sqmuxa_i_TMR_0(main_basesoc_serial_tx_rs232phytx_next_value1_1_sqmuxa_i_TMR_0),
    .main_basesoc_serial_tx_rs232phytx_next_value1_1_sqmuxa_i_TMR_1(main_basesoc_serial_tx_rs232phytx_next_value1_1_sqmuxa_i_TMR_1),
    .main_basesoc_serial_tx_rs232phytx_next_value1_1_sqmuxa_i_TMR_2(main_basesoc_serial_tx_rs232phytx_next_value1_1_sqmuxa_i_TMR_2),
    .main_basesoc_timer_en_storage_TMR_0(main_basesoc_timer_en_storage_TMR_0),
    .main_basesoc_timer_en_storage_TMR_1(main_basesoc_timer_en_storage_TMR_1),
    .main_basesoc_timer_en_storage_TMR_2(main_basesoc_timer_en_storage_TMR_2),
    .main_basesoc_timer_enable_storage_TMR_0(main_basesoc_timer_enable_storage_TMR_0),
    .main_basesoc_timer_enable_storage_TMR_1(main_basesoc_timer_enable_storage_TMR_1),
    .main_basesoc_timer_enable_storage_TMR_2(main_basesoc_timer_enable_storage_TMR_2),
    .main_basesoc_timer_pending_r_0_sqmuxa_1z_TMR_0(main_basesoc_timer_pending_r_0_sqmuxa_TMR_0),
    .main_basesoc_timer_pending_r_0_sqmuxa_1z_TMR_1(main_basesoc_timer_pending_r_0_sqmuxa_TMR_1),
    .main_basesoc_timer_pending_r_0_sqmuxa_1z_TMR_2(main_basesoc_timer_pending_r_0_sqmuxa_TMR_2),
    .main_basesoc_timer_pending_r_TMR_0(main_basesoc_timer_pending_r_TMR_0),
    .main_basesoc_timer_pending_r_TMR_1(main_basesoc_timer_pending_r_TMR_1),
    .main_basesoc_timer_pending_r_TMR_2(main_basesoc_timer_pending_r_TMR_2),
    .main_basesoc_timer_pending_re_TMR_0(main_basesoc_timer_pending_re_TMR_0),
    .main_basesoc_timer_pending_re_TMR_1(main_basesoc_timer_pending_re_TMR_1),
    .main_basesoc_timer_pending_re_TMR_2(main_basesoc_timer_pending_re_TMR_2),
    .main_basesoc_timer_reload_storage_TMR_0(main_basesoc_timer_reload_storage_TMR_0),
    .main_basesoc_timer_reload_storage_TMR_1(main_basesoc_timer_reload_storage_TMR_1),
    .main_basesoc_timer_reload_storage_TMR_2(main_basesoc_timer_reload_storage_TMR_2),
    .main_basesoc_timer_update_value_storage_0_sqmuxa_1z_TMR_0(main_basesoc_timer_update_value_storage_0_sqmuxa_TMR_0),
    .main_basesoc_timer_update_value_storage_0_sqmuxa_1z_TMR_1(main_basesoc_timer_update_value_storage_0_sqmuxa_TMR_1),
    .main_basesoc_timer_update_value_storage_0_sqmuxa_1z_TMR_2(main_basesoc_timer_update_value_storage_0_sqmuxa_TMR_2),
    .main_basesoc_timer_update_value_storage_TMR_0(main_basesoc_timer_update_value_storage_TMR_0),
    .main_basesoc_timer_update_value_storage_TMR_1(main_basesoc_timer_update_value_storage_TMR_1),
    .main_basesoc_timer_update_value_storage_TMR_2(main_basesoc_timer_update_value_storage_TMR_2),
    .main_basesoc_timer_value_7_0_0_TMR_0(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_0_0_TMR_0 ),
    .main_basesoc_timer_value_7_0_0_TMR_1(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_0_0_TMR_1 ),
    .main_basesoc_timer_value_7_0_0_TMR_2(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_0_0_TMR_2 ),
    .main_basesoc_timer_value_7_1_TMR_0(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 ),
    .main_basesoc_timer_value_7_1_TMR_1(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 ),
    .main_basesoc_timer_value_7_1_TMR_2(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 ),
    .main_basesoc_timer_value_7_TMR_0(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_0 ),
    .main_basesoc_timer_value_7_TMR_1(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_1 ),
    .main_basesoc_timer_value_7_TMR_2(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_2 ),
    .main_basesoc_timer_value_status_TMR_0(main_basesoc_timer_value_status_TMR_0),
    .main_basesoc_timer_value_status_TMR_1(main_basesoc_timer_value_status_TMR_1),
    .main_basesoc_timer_value_status_TMR_2(main_basesoc_timer_value_status_TMR_2),
    .main_basesoc_timer_zero_pending_TMR_0(main_basesoc_timer_zero_pending_TMR_0),
    .main_basesoc_timer_zero_pending_TMR_1(main_basesoc_timer_zero_pending_TMR_1),
    .main_basesoc_timer_zero_pending_TMR_2(main_basesoc_timer_zero_pending_TMR_2),
    .main_basesoc_timer_zero_trigger_TMR_0(main_basesoc_timer_zero_trigger_TMR_0),
    .main_basesoc_timer_zero_trigger_TMR_1(main_basesoc_timer_zero_trigger_TMR_1),
    .main_basesoc_timer_zero_trigger_TMR_2(main_basesoc_timer_zero_trigger_TMR_2),
    .main_basesoc_timer_zero_trigger_d_TMR_0(main_basesoc_timer_zero_trigger_d_TMR_0),
    .main_basesoc_timer_zero_trigger_d_TMR_1(main_basesoc_timer_zero_trigger_d_TMR_1),
    .main_basesoc_timer_zero_trigger_d_TMR_2(main_basesoc_timer_zero_trigger_d_TMR_2),
    .main_basesoc_tx_count_TMR_0(main_basesoc_tx_count_TMR_0),
    .main_basesoc_tx_count_TMR_1(main_basesoc_tx_count_TMR_1),
    .main_basesoc_tx_count_TMR_2(main_basesoc_tx_count_TMR_2),
    .main_basesoc_tx_count_rs232phytx_next_value0_TMR_0(main_basesoc_tx_count_rs232phytx_next_value0_TMR_0),
    .main_basesoc_tx_count_rs232phytx_next_value0_TMR_1(main_basesoc_tx_count_rs232phytx_next_value0_TMR_1),
    .main_basesoc_tx_count_rs232phytx_next_value0_TMR_2(main_basesoc_tx_count_rs232phytx_next_value0_TMR_2),
    .main_basesoc_tx_data_TMR_0(main_basesoc_tx_data_TMR_0),
    .main_basesoc_tx_data_TMR_1(main_basesoc_tx_data_TMR_1),
    .main_basesoc_tx_data_TMR_2(main_basesoc_tx_data_TMR_2),
    .main_basesoc_tx_data_rs232phytx_next_value2_0_sqmuxa_TMR_0(main_basesoc_tx_data_rs232phytx_next_value2_0_sqmuxa_TMR_0),
    .main_basesoc_tx_data_rs232phytx_next_value2_0_sqmuxa_TMR_1(main_basesoc_tx_data_rs232phytx_next_value2_0_sqmuxa_TMR_1),
    .main_basesoc_tx_data_rs232phytx_next_value2_0_sqmuxa_TMR_2(main_basesoc_tx_data_rs232phytx_next_value2_0_sqmuxa_TMR_2),
    .main_basesoc_tx_data_rs232phytx_next_value2_TMR_0(main_basesoc_tx_data_rs232phytx_next_value2_TMR_0),
    .main_basesoc_tx_data_rs232phytx_next_value2_TMR_1(main_basesoc_tx_data_rs232phytx_next_value2_TMR_1),
    .main_basesoc_tx_data_rs232phytx_next_value2_TMR_2(main_basesoc_tx_data_rs232phytx_next_value2_TMR_2),
    .main_basesoc_tx_data_rs232phytx_next_value_ce2_1_TMR_0(main_basesoc_tx_data_rs232phytx_next_value_ce2_1_TMR_0),
    .main_basesoc_tx_data_rs232phytx_next_value_ce2_1_TMR_1(main_basesoc_tx_data_rs232phytx_next_value_ce2_1_TMR_1),
    .main_basesoc_tx_data_rs232phytx_next_value_ce2_1_TMR_2(main_basesoc_tx_data_rs232phytx_next_value_ce2_1_TMR_2),
    .main_basesoc_tx_tick_0_TMR_0(main_basesoc_tx_tick_0_TMR_0),
    .main_basesoc_tx_tick_0_TMR_1(main_basesoc_tx_tick_0_TMR_1),
    .main_basesoc_tx_tick_0_TMR_2(main_basesoc_tx_tick_0_TMR_2),
    .main_basesoc_tx_tick_TMR_0(main_basesoc_tx_tick_TMR_0),
    .main_basesoc_tx_tick_TMR_1(main_basesoc_tx_tick_TMR_1),
    .main_basesoc_tx_tick_TMR_2(main_basesoc_tx_tick_TMR_2),
    .main_basesoc_uart_enable_storage_TMR_0(main_basesoc_uart_enable_storage_TMR_0),
    .main_basesoc_uart_enable_storage_TMR_1(main_basesoc_uart_enable_storage_TMR_1),
    .main_basesoc_uart_enable_storage_TMR_2(main_basesoc_uart_enable_storage_TMR_2),
    .main_basesoc_uart_pending_r_0_sqmuxa_1z_TMR_0(main_basesoc_uart_pending_r_0_sqmuxa_TMR_0),
    .main_basesoc_uart_pending_r_0_sqmuxa_1z_TMR_1(main_basesoc_uart_pending_r_0_sqmuxa_TMR_1),
    .main_basesoc_uart_pending_r_0_sqmuxa_1z_TMR_2(main_basesoc_uart_pending_r_0_sqmuxa_TMR_2),
    .main_basesoc_uart_pending_r_TMR_0(main_basesoc_uart_pending_r_TMR_0),
    .main_basesoc_uart_pending_r_TMR_1(main_basesoc_uart_pending_r_TMR_1),
    .main_basesoc_uart_pending_r_TMR_2(main_basesoc_uart_pending_r_TMR_2),
    .main_basesoc_uart_pending_re_TMR_0(main_basesoc_uart_pending_re_TMR_0),
    .main_basesoc_uart_pending_re_TMR_1(main_basesoc_uart_pending_re_TMR_1),
    .main_basesoc_uart_pending_re_TMR_2(main_basesoc_uart_pending_re_TMR_2),
    .main_basesoc_uart_rx_fifo_readable_TMR_0(main_basesoc_uart_rx_fifo_readable_TMR_0),
    .main_basesoc_uart_rx_fifo_readable_TMR_1(main_basesoc_uart_rx_fifo_readable_TMR_1),
    .main_basesoc_uart_rx_fifo_readable_TMR_2(main_basesoc_uart_rx_fifo_readable_TMR_2),
    .main_basesoc_uart_rx_fifo_syncfifo_re_TMR_0(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_0),
    .main_basesoc_uart_rx_fifo_syncfifo_re_TMR_1(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_1),
    .main_basesoc_uart_rx_fifo_syncfifo_re_TMR_2(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_2),
    .main_basesoc_uart_rx_fifo_wrport_we_TMR_0(main_basesoc_uart_rx_fifo_wrport_we_TMR_0),
    .main_basesoc_uart_rx_fifo_wrport_we_TMR_1(main_basesoc_uart_rx_fifo_wrport_we_TMR_1),
    .main_basesoc_uart_rx_fifo_wrport_we_TMR_2(main_basesoc_uart_rx_fifo_wrport_we_TMR_2),
    .main_basesoc_uart_rx_pending_TMR_0(main_basesoc_uart_rx_pending_TMR_0),
    .main_basesoc_uart_rx_pending_TMR_1(main_basesoc_uart_rx_pending_TMR_1),
    .main_basesoc_uart_rx_pending_TMR_2(main_basesoc_uart_rx_pending_TMR_2),
    .main_basesoc_uart_rx_trigger_d_TMR_0(main_basesoc_uart_rx_trigger_d_TMR_0),
    .main_basesoc_uart_rx_trigger_d_TMR_1(main_basesoc_uart_rx_trigger_d_TMR_1),
    .main_basesoc_uart_rx_trigger_d_TMR_2(main_basesoc_uart_rx_trigger_d_TMR_2),
    .main_basesoc_uart_tx_fifo_level0_0_mod_RNIG0F3_0_TMR_0(main_basesoc_uart_tx_fifo_level0_0_mod_RNIG0F3_TMR_0),
    .main_basesoc_uart_tx_fifo_level0_0_mod_RNIG0F3_0_TMR_1(main_basesoc_uart_tx_fifo_level0_0_mod_RNIG0F3_TMR_1),
    .main_basesoc_uart_tx_fifo_level0_0_mod_RNIG0F3_0_TMR_2(main_basesoc_uart_tx_fifo_level0_0_mod_RNIG0F3_TMR_2),
    .main_basesoc_uart_tx_fifo_readable_TMR_0(main_basesoc_uart_tx_fifo_readable_TMR_0),
    .main_basesoc_uart_tx_fifo_readable_TMR_1(main_basesoc_uart_tx_fifo_readable_TMR_1),
    .main_basesoc_uart_tx_fifo_readable_TMR_2(main_basesoc_uart_tx_fifo_readable_TMR_2),
    .main_basesoc_uart_tx_fifo_syncfifo_re_TMR_0(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_0),
    .main_basesoc_uart_tx_fifo_syncfifo_re_TMR_1(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_1),
    .main_basesoc_uart_tx_fifo_syncfifo_re_TMR_2(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_2),
    .main_basesoc_uart_tx_fifo_wrport_we_TMR_0(main_basesoc_uart_tx_fifo_wrport_we_TMR_0),
    .main_basesoc_uart_tx_fifo_wrport_we_TMR_1(main_basesoc_uart_tx_fifo_wrport_we_TMR_1),
    .main_basesoc_uart_tx_fifo_wrport_we_TMR_2(main_basesoc_uart_tx_fifo_wrport_we_TMR_2),
    .main_basesoc_uart_tx_pending_TMR_0(main_basesoc_uart_tx_pending_TMR_0),
    .main_basesoc_uart_tx_pending_TMR_1(main_basesoc_uart_tx_pending_TMR_1),
    .main_basesoc_uart_tx_pending_TMR_2(main_basesoc_uart_tx_pending_TMR_2),
    .main_basesoc_uart_tx_trigger_d_TMR_0(main_basesoc_uart_tx_trigger_d_TMR_0),
    .main_basesoc_uart_tx_trigger_d_TMR_1(main_basesoc_uart_tx_trigger_d_TMR_1),
    .main_basesoc_uart_tx_trigger_d_TMR_2(main_basesoc_uart_tx_trigger_d_TMR_2),
    .main_bus_ack_TMR_0(main_bus_ack_TMR_0),
    .main_bus_ack_TMR_1(main_bus_ack_TMR_1),
    .main_bus_ack_TMR_2(main_bus_ack_TMR_2),
    .main_bus_ack_r_0_a2_TMR_0(main_bus_ack_r_0_a2_TMR_0),
    .main_bus_ack_r_0_a2_TMR_1(main_bus_ack_r_0_a2_TMR_1),
    .main_bus_ack_r_0_a2_TMR_2(main_bus_ack_r_0_a2_TMR_2),
    .main_chaser_TMR_0(main_chaser_TMR_0),
    .main_chaser_TMR_1(main_chaser_TMR_1),
    .main_chaser_TMR_2(main_chaser_TMR_2),
    .main_cs06_TMR_0(main_cs06_TMR_0),
    .main_cs06_TMR_1(main_cs06_TMR_1),
    .main_cs06_TMR_2(main_cs06_TMR_2),
    .main_dataout0(main_dataout0),
    .main_dataout1(main_dataout1),
    .main_m1_e_0_1_TMR_0(\VexRiscv.main_m1_e_0_1_TMR_0 ),
    .main_m1_e_0_1_TMR_1(\VexRiscv.main_m1_e_0_1_TMR_1 ),
    .main_m1_e_0_1_TMR_2(\VexRiscv.main_m1_e_0_1_TMR_2 ),
    .main_mode_TMR_0(main_mode_TMR_0),
    .main_mode_TMR_1(main_mode_TMR_1),
    .main_mode_TMR_2(main_mode_TMR_2),
    .main_storage_0_sqmuxa_TMR_0(main_storage_0_sqmuxa_TMR_0),
    .main_storage_0_sqmuxa_TMR_1(main_storage_0_sqmuxa_TMR_1),
    .main_storage_0_sqmuxa_TMR_2(main_storage_0_sqmuxa_TMR_2),
    .main_storage_TMR_0(main_storage_TMR_0),
    .main_storage_TMR_1(main_storage_TMR_1),
    .main_storage_TMR_2(main_storage_TMR_2),
    .main_wren0_TMR_0(main_wren0_TMR_0),
    .main_wren0_TMR_1(main_wren0_TMR_1),
    .main_wren0_TMR_2(main_wren0_TMR_2),
    .main_wren1_TMR_0(main_wren1_TMR_0),
    .main_wren1_TMR_1(main_wren1_TMR_1),
    .main_wren1_TMR_2(main_wren1_TMR_2),
    .rom_dat0(rom_dat0),
    .serial_tx_4_TMR_0(serial_tx_4_TMR_0),
    .serial_tx_4_TMR_1(serial_tx_4_TMR_1),
    .serial_tx_4_TMR_2(serial_tx_4_TMR_2),
    .storage_1_dat1_TMR_0(storage_1_dat1_TMR_0[1:0]),
    .storage_1_dat1_TMR_1(storage_1_dat1_TMR_1[1:0]),
    .storage_1_dat1_TMR_2(storage_1_dat1_TMR_2[1:0]),
    .storage_dat1_TMR_0(storage_dat1_TMR_0),
    .storage_dat1_TMR_1(storage_dat1_TMR_1),
    .storage_dat1_TMR_2(storage_dat1_TMR_2),
    .sys_clk_0(sys_clk),
    .sys_rst_TMR_0(sys_rst_TMR_0),
    .sys_rst_TMR_1(sys_rst_TMR_1),
    .sys_rst_TMR_2(sys_rst_TMR_2),
    .un1_main_basesoc_bus_errors_1_0_TMR_0(un1_main_basesoc_bus_errors_1_0_TMR_0),
    .un1_main_basesoc_bus_errors_1_0_TMR_1(un1_main_basesoc_bus_errors_1_0_TMR_1),
    .un1_main_basesoc_bus_errors_1_0_TMR_2(un1_main_basesoc_bus_errors_1_0_TMR_2),
    .un1_main_basesoc_serial_tx_rs232phytx_next_value112_i_0_TMR_0(un1_main_basesoc_serial_tx_rs232phytx_next_value112_i_TMR_0),
    .un1_main_basesoc_serial_tx_rs232phytx_next_value112_i_0_TMR_1(un1_main_basesoc_serial_tx_rs232phytx_next_value112_i_TMR_1),
    .un1_main_basesoc_serial_tx_rs232phytx_next_value112_i_0_TMR_2(un1_main_basesoc_serial_tx_rs232phytx_next_value112_i_TMR_2),
    .un1_main_basesoc_uart_rx_fifo_level0_0_TMR_0(un1_main_basesoc_uart_rx_fifo_level0_0_TMR_0),
    .un1_main_basesoc_uart_rx_fifo_level0_0_TMR_1(un1_main_basesoc_uart_rx_fifo_level0_0_TMR_1),
    .un1_main_basesoc_uart_rx_fifo_level0_0_TMR_2(un1_main_basesoc_uart_rx_fifo_level0_0_TMR_2),
    .un1_main_basesoc_uart_rx_fifo_level0_TMR_0(un1_main_basesoc_uart_rx_fifo_level0_scalar_TMR_0),
    .un1_main_basesoc_uart_rx_fifo_level0_TMR_1(un1_main_basesoc_uart_rx_fifo_level0_scalar_TMR_1),
    .un1_main_basesoc_uart_rx_fifo_level0_TMR_2(un1_main_basesoc_uart_rx_fifo_level0_scalar_TMR_2),
    .un1_main_basesoc_uart_tx_fifo_level0_0_TMR_0(un1_main_basesoc_uart_tx_fifo_level0_0_TMR_0),
    .un1_main_basesoc_uart_tx_fifo_level0_0_TMR_1(un1_main_basesoc_uart_tx_fifo_level0_0_TMR_1),
    .un1_main_basesoc_uart_tx_fifo_level0_0_TMR_2(un1_main_basesoc_uart_tx_fifo_level0_0_TMR_2),
    .un1_main_basesoc_uart_tx_fifo_level0_0_d0_TMR_0(un1_main_basesoc_uart_tx_fifo_level0_TMR_0[0]),
    .un1_main_basesoc_uart_tx_fifo_level0_0_d0_TMR_1(un1_main_basesoc_uart_tx_fifo_level0_TMR_1[0]),
    .un1_main_basesoc_uart_tx_fifo_level0_0_d0_TMR_2(un1_main_basesoc_uart_tx_fifo_level0_TMR_2[0]),
    .un1_main_basesoc_uart_tx_fifo_level0_1z_TMR_0(un1_main_basesoc_uart_tx_fifo_level0_scalar_TMR_0),
    .un1_main_basesoc_uart_tx_fifo_level0_1z_TMR_1(un1_main_basesoc_uart_tx_fifo_level0_scalar_TMR_1),
    .un1_main_basesoc_uart_tx_fifo_level0_1z_TMR_2(un1_main_basesoc_uart_tx_fifo_level0_scalar_TMR_2),
    .un1_main_basesoc_uart_tx_fifo_produce_axbxc3_m6_e_3_TMR_0(un1_main_basesoc_uart_tx_fifo_produce_axbxc3_m6_e_3_TMR_0),
    .un1_main_basesoc_uart_tx_fifo_produce_axbxc3_m6_e_3_TMR_1(un1_main_basesoc_uart_tx_fifo_produce_axbxc3_m6_e_3_TMR_1),
    .un1_main_basesoc_uart_tx_fifo_produce_axbxc3_m6_e_3_TMR_2(un1_main_basesoc_uart_tx_fifo_produce_axbxc3_m6_e_3_TMR_2),
    .un3_main_basesoc_uart_tx_fifo_syncfifo_writable_i_TMR_0(un3_main_basesoc_uart_tx_fifo_syncfifo_writable_i_TMR_0),
    .un3_main_basesoc_uart_tx_fifo_syncfifo_writable_i_TMR_1(un3_main_basesoc_uart_tx_fifo_syncfifo_writable_i_TMR_1),
    .un3_main_basesoc_uart_tx_fifo_syncfifo_writable_i_TMR_2(un3_main_basesoc_uart_tx_fifo_syncfifo_writable_i_TMR_2),
    .un5_main_basesoc_rx_phase_cry_31_TMR_0(un5_main_basesoc_rx_phase_cry_31_TMR_0),
    .un5_main_basesoc_rx_phase_cry_31_TMR_1(un5_main_basesoc_rx_phase_cry_31_TMR_1),
    .un5_main_basesoc_rx_phase_cry_31_TMR_2(un5_main_basesoc_rx_phase_cry_31_TMR_2),
    .un5_main_basesoc_tx_phase_cry_31_TMR_0(un5_main_basesoc_tx_phase_cry_31_TMR_0),
    .un5_main_basesoc_tx_phase_cry_31_TMR_1(un5_main_basesoc_tx_phase_cry_31_TMR_1),
    .un5_main_basesoc_tx_phase_cry_31_TMR_2(un5_main_basesoc_tx_phase_cry_31_TMR_2),
    .user_led0_c_TMR_0(user_led0_c_TMR_0),
    .user_led0_c_TMR_1(user_led0_c_TMR_1),
    .user_led0_c_TMR_2(user_led0_c_TMR_2),
    .user_led10_c_TMR_0(user_led10_c_TMR_0),
    .user_led10_c_TMR_1(user_led10_c_TMR_1),
    .user_led10_c_TMR_2(user_led10_c_TMR_2),
    .user_led11_c_TMR_0(user_led11_c_TMR_0),
    .user_led11_c_TMR_1(user_led11_c_TMR_1),
    .user_led11_c_TMR_2(user_led11_c_TMR_2),
    .user_led12_c_TMR_0(user_led12_c_TMR_0),
    .user_led12_c_TMR_1(user_led12_c_TMR_1),
    .user_led12_c_TMR_2(user_led12_c_TMR_2),
    .user_led13_c_TMR_0(user_led13_c_TMR_0),
    .user_led13_c_TMR_1(user_led13_c_TMR_1),
    .user_led13_c_TMR_2(user_led13_c_TMR_2),
    .user_led1_c_TMR_0(user_led1_c_TMR_0),
    .user_led1_c_TMR_1(user_led1_c_TMR_1),
    .user_led1_c_TMR_2(user_led1_c_TMR_2),
    .user_led2_c_TMR_0(user_led2_c_TMR_0),
    .user_led2_c_TMR_1(user_led2_c_TMR_1),
    .user_led2_c_TMR_2(user_led2_c_TMR_2),
    .user_led3_c_TMR_0(user_led3_c_TMR_0),
    .user_led3_c_TMR_1(user_led3_c_TMR_1),
    .user_led3_c_TMR_2(user_led3_c_TMR_2),
    .user_led4_c_TMR_0(user_led4_c_TMR_0),
    .user_led4_c_TMR_1(user_led4_c_TMR_1),
    .user_led4_c_TMR_2(user_led4_c_TMR_2),
    .user_led5_c_TMR_0(user_led5_c_TMR_0),
    .user_led5_c_TMR_1(user_led5_c_TMR_1),
    .user_led5_c_TMR_2(user_led5_c_TMR_2),
    .user_led6_c_TMR_0(user_led6_c_TMR_0),
    .user_led6_c_TMR_1(user_led6_c_TMR_1),
    .user_led6_c_TMR_2(user_led6_c_TMR_2),
    .user_led7_c_TMR_0(user_led7_c_TMR_0),
    .user_led7_c_TMR_1(user_led7_c_TMR_1),
    .user_led7_c_TMR_2(user_led7_c_TMR_2),
    .user_led8_c_TMR_0(user_led8_c_TMR_0),
    .user_led8_c_TMR_1(user_led8_c_TMR_1),
    .user_led8_c_TMR_2(user_led8_c_TMR_2),
    .user_led9_c_TMR_0(user_led9_c_TMR_0),
    .user_led9_c_TMR_1(user_led9_c_TMR_1),
    .user_led9_c_TMR_2(user_led9_c_TMR_2)
  );
  LUT4 builder_array_muxed0_0_RED_VOTER (
    .A(builder_array_muxed0_TMR_0[0]),
    .B(builder_array_muxed0_TMR_1[0]),
    .C(builder_array_muxed0_TMR_2[0]),
    .D(1'h0),
    .Z(builder_array_muxed0_0_RED_VOTER_wire)
  );
  defparam builder_array_muxed0_0_RED_VOTER.INIT = "0xFCC0";
  LUT4 builder_array_muxed0_10_RED_VOTER (
    .A(builder_array_muxed0_TMR_0[10]),
    .B(builder_array_muxed0_TMR_1[10]),
    .C(builder_array_muxed0_TMR_2[10]),
    .D(1'h0),
    .Z(builder_array_muxed0_10_RED_VOTER_wire)
  );
  defparam builder_array_muxed0_10_RED_VOTER.INIT = "0xFCC0";
  LUT4 builder_array_muxed0_11_RED_VOTER (
    .A(builder_array_muxed0_TMR_0[11]),
    .B(builder_array_muxed0_TMR_1[11]),
    .C(builder_array_muxed0_TMR_2[11]),
    .D(1'h0),
    .Z(builder_array_muxed0_11_RED_VOTER_wire)
  );
  defparam builder_array_muxed0_11_RED_VOTER.INIT = "0xFCC0";
  LUT4 builder_array_muxed0_12_RED_VOTER (
    .A(builder_array_muxed0_TMR_0[12]),
    .B(builder_array_muxed0_TMR_1[12]),
    .C(builder_array_muxed0_TMR_2[12]),
    .D(1'h0),
    .Z(builder_array_muxed0_12_RED_VOTER_wire)
  );
  defparam builder_array_muxed0_12_RED_VOTER.INIT = "0xFCC0";
  LUT4 builder_array_muxed0_13_RED_VOTER (
    .A(builder_array_muxed0_TMR_0[13]),
    .B(builder_array_muxed0_TMR_1[13]),
    .C(builder_array_muxed0_TMR_2[13]),
    .D(1'h0),
    .Z(builder_array_muxed0_13_RED_VOTER_wire)
  );
  defparam builder_array_muxed0_13_RED_VOTER.INIT = "0xFCC0";
  LUT4 builder_array_muxed0_1_RED_VOTER (
    .A(builder_array_muxed0_TMR_0[1]),
    .B(builder_array_muxed0_TMR_1[1]),
    .C(builder_array_muxed0_TMR_2[1]),
    .D(1'h0),
    .Z(builder_array_muxed0_1_RED_VOTER_wire)
  );
  defparam builder_array_muxed0_1_RED_VOTER.INIT = "0xFCC0";
  LUT4 builder_array_muxed0_2_RED_VOTER (
    .A(builder_array_muxed0_TMR_0[2]),
    .B(builder_array_muxed0_TMR_1[2]),
    .C(builder_array_muxed0_TMR_2[2]),
    .D(1'h0),
    .Z(builder_array_muxed0_2_RED_VOTER_wire)
  );
  defparam builder_array_muxed0_2_RED_VOTER.INIT = "0xFCC0";
  LUT4 builder_array_muxed0_4_RED_VOTER (
    .A(builder_array_muxed0_TMR_0[4]),
    .B(builder_array_muxed0_TMR_1[4]),
    .C(builder_array_muxed0_TMR_2[4]),
    .D(1'h0),
    .Z(builder_array_muxed0_4_RED_VOTER_wire)
  );
  defparam builder_array_muxed0_4_RED_VOTER.INIT = "0xFCC0";
  LUT4 builder_array_muxed0_5_RED_VOTER (
    .A(builder_array_muxed0_TMR_0[5]),
    .B(builder_array_muxed0_TMR_1[5]),
    .C(builder_array_muxed0_TMR_2[5]),
    .D(1'h0),
    .Z(builder_array_muxed0_5_RED_VOTER_wire)
  );
  defparam builder_array_muxed0_5_RED_VOTER.INIT = "0xFCC0";
  LUT4 builder_array_muxed0_6_RED_VOTER (
    .A(builder_array_muxed0_TMR_0[6]),
    .B(builder_array_muxed0_TMR_1[6]),
    .C(builder_array_muxed0_TMR_2[6]),
    .D(1'h0),
    .Z(builder_array_muxed0_6_RED_VOTER_wire)
  );
  defparam builder_array_muxed0_6_RED_VOTER.INIT = "0xFCC0";
  LUT4 builder_array_muxed0_7_RED_VOTER (
    .A(builder_array_muxed0_TMR_0[7]),
    .B(builder_array_muxed0_TMR_1[7]),
    .C(builder_array_muxed0_TMR_2[7]),
    .D(1'h0),
    .Z(builder_array_muxed0_7_RED_VOTER_wire)
  );
  defparam builder_array_muxed0_7_RED_VOTER.INIT = "0xFCC0";
  LUT4 builder_array_muxed0_8_RED_VOTER (
    .A(builder_array_muxed0_TMR_0[8]),
    .B(builder_array_muxed0_TMR_1[8]),
    .C(builder_array_muxed0_TMR_2[8]),
    .D(1'h0),
    .Z(builder_array_muxed0_8_RED_VOTER_wire)
  );
  defparam builder_array_muxed0_8_RED_VOTER.INIT = "0xFCC0";
  LUT4 builder_array_muxed0_9_RED_VOTER (
    .A(builder_array_muxed0_TMR_0[9]),
    .B(builder_array_muxed0_TMR_1[9]),
    .C(builder_array_muxed0_TMR_2[9]),
    .D(1'h0),
    .Z(builder_array_muxed0_9_RED_VOTER_wire)
  );
  defparam builder_array_muxed0_9_RED_VOTER.INIT = "0xFCC0";
  LUT4 builder_array_muxed1_0_RED_VOTER (
    .A(builder_array_muxed1_TMR_0[0]),
    .B(builder_array_muxed1_TMR_1[0]),
    .C(builder_array_muxed1_TMR_2[0]),
    .D(1'h0),
    .Z(builder_array_muxed1_0_RED_VOTER_wire)
  );
  defparam builder_array_muxed1_0_RED_VOTER.INIT = "0xFCC0";
  LUT4 builder_array_muxed1_10_RED_VOTER (
    .A(builder_array_muxed1_TMR_0[10]),
    .B(builder_array_muxed1_TMR_1[10]),
    .C(builder_array_muxed1_TMR_2[10]),
    .D(1'h0),
    .Z(builder_array_muxed1_10_RED_VOTER_wire)
  );
  defparam builder_array_muxed1_10_RED_VOTER.INIT = "0xFCC0";
  LUT4 builder_array_muxed1_11_RED_VOTER (
    .A(builder_array_muxed1_TMR_0[11]),
    .B(builder_array_muxed1_TMR_1[11]),
    .C(builder_array_muxed1_TMR_2[11]),
    .D(1'h0),
    .Z(builder_array_muxed1_11_RED_VOTER_wire)
  );
  defparam builder_array_muxed1_11_RED_VOTER.INIT = "0xFCC0";
  LUT4 builder_array_muxed1_12_RED_VOTER (
    .A(builder_array_muxed1_TMR_0[12]),
    .B(builder_array_muxed1_TMR_1[12]),
    .C(builder_array_muxed1_TMR_2[12]),
    .D(1'h0),
    .Z(builder_array_muxed1_12_RED_VOTER_wire)
  );
  defparam builder_array_muxed1_12_RED_VOTER.INIT = "0xFCC0";
  LUT4 builder_array_muxed1_13_RED_VOTER (
    .A(builder_array_muxed1_TMR_0[13]),
    .B(builder_array_muxed1_TMR_1[13]),
    .C(builder_array_muxed1_TMR_2[13]),
    .D(1'h0),
    .Z(builder_array_muxed1_13_RED_VOTER_wire)
  );
  defparam builder_array_muxed1_13_RED_VOTER.INIT = "0xFCC0";
  LUT4 builder_array_muxed1_14_RED_VOTER (
    .A(builder_array_muxed1_TMR_0[14]),
    .B(builder_array_muxed1_TMR_1[14]),
    .C(builder_array_muxed1_TMR_2[14]),
    .D(1'h0),
    .Z(builder_array_muxed1_14_RED_VOTER_wire)
  );
  defparam builder_array_muxed1_14_RED_VOTER.INIT = "0xFCC0";
  LUT4 builder_array_muxed1_15_RED_VOTER (
    .A(builder_array_muxed1_TMR_0[15]),
    .B(builder_array_muxed1_TMR_1[15]),
    .C(builder_array_muxed1_TMR_2[15]),
    .D(1'h0),
    .Z(builder_array_muxed1_15_RED_VOTER_wire)
  );
  defparam builder_array_muxed1_15_RED_VOTER.INIT = "0xFCC0";
  LUT4 builder_array_muxed1_16_RED_VOTER (
    .A(builder_array_muxed1_TMR_0[16]),
    .B(builder_array_muxed1_TMR_1[16]),
    .C(builder_array_muxed1_TMR_2[16]),
    .D(1'h0),
    .Z(builder_array_muxed1_16_RED_VOTER_wire)
  );
  defparam builder_array_muxed1_16_RED_VOTER.INIT = "0xFCC0";
  LUT4 builder_array_muxed1_17_RED_VOTER (
    .A(builder_array_muxed1_TMR_0[17]),
    .B(builder_array_muxed1_TMR_1[17]),
    .C(builder_array_muxed1_TMR_2[17]),
    .D(1'h0),
    .Z(builder_array_muxed1_17_RED_VOTER_wire)
  );
  defparam builder_array_muxed1_17_RED_VOTER.INIT = "0xFCC0";
  LUT4 builder_array_muxed1_18_RED_VOTER (
    .A(builder_array_muxed1_TMR_0[18]),
    .B(builder_array_muxed1_TMR_1[18]),
    .C(builder_array_muxed1_TMR_2[18]),
    .D(1'h0),
    .Z(builder_array_muxed1_18_RED_VOTER_wire)
  );
  defparam builder_array_muxed1_18_RED_VOTER.INIT = "0xFCC0";
  LUT4 builder_array_muxed1_19_RED_VOTER (
    .A(builder_array_muxed1_TMR_0[19]),
    .B(builder_array_muxed1_TMR_1[19]),
    .C(builder_array_muxed1_TMR_2[19]),
    .D(1'h0),
    .Z(builder_array_muxed1_19_RED_VOTER_wire)
  );
  defparam builder_array_muxed1_19_RED_VOTER.INIT = "0xFCC0";
  LUT4 builder_array_muxed1_1_RED_VOTER (
    .A(builder_array_muxed1_TMR_0[1]),
    .B(builder_array_muxed1_TMR_1[1]),
    .C(builder_array_muxed1_TMR_2[1]),
    .D(1'h0),
    .Z(builder_array_muxed1_1_RED_VOTER_wire)
  );
  defparam builder_array_muxed1_1_RED_VOTER.INIT = "0xFCC0";
  LUT4 builder_array_muxed1_20_RED_VOTER (
    .A(builder_array_muxed1_TMR_0[20]),
    .B(builder_array_muxed1_TMR_1[20]),
    .C(builder_array_muxed1_TMR_2[20]),
    .D(1'h0),
    .Z(builder_array_muxed1_20_RED_VOTER_wire)
  );
  defparam builder_array_muxed1_20_RED_VOTER.INIT = "0xFCC0";
  LUT4 builder_array_muxed1_21_RED_VOTER (
    .A(builder_array_muxed1_TMR_0[21]),
    .B(builder_array_muxed1_TMR_1[21]),
    .C(builder_array_muxed1_TMR_2[21]),
    .D(1'h0),
    .Z(builder_array_muxed1_21_RED_VOTER_wire)
  );
  defparam builder_array_muxed1_21_RED_VOTER.INIT = "0xFCC0";
  LUT4 builder_array_muxed1_22_RED_VOTER (
    .A(builder_array_muxed1_TMR_0[22]),
    .B(builder_array_muxed1_TMR_1[22]),
    .C(builder_array_muxed1_TMR_2[22]),
    .D(1'h0),
    .Z(builder_array_muxed1_22_RED_VOTER_wire)
  );
  defparam builder_array_muxed1_22_RED_VOTER.INIT = "0xFCC0";
  LUT4 builder_array_muxed1_23_RED_VOTER (
    .A(builder_array_muxed1_TMR_0[23]),
    .B(builder_array_muxed1_TMR_1[23]),
    .C(builder_array_muxed1_TMR_2[23]),
    .D(1'h0),
    .Z(builder_array_muxed1_23_RED_VOTER_wire)
  );
  defparam builder_array_muxed1_23_RED_VOTER.INIT = "0xFCC0";
  LUT4 builder_array_muxed1_24_RED_VOTER (
    .A(builder_array_muxed1_TMR_0[24]),
    .B(builder_array_muxed1_TMR_1[24]),
    .C(builder_array_muxed1_TMR_2[24]),
    .D(1'h0),
    .Z(builder_array_muxed1_24_RED_VOTER_wire)
  );
  defparam builder_array_muxed1_24_RED_VOTER.INIT = "0xFCC0";
  LUT4 builder_array_muxed1_25_RED_VOTER (
    .A(builder_array_muxed1_TMR_0[25]),
    .B(builder_array_muxed1_TMR_1[25]),
    .C(builder_array_muxed1_TMR_2[25]),
    .D(1'h0),
    .Z(builder_array_muxed1_25_RED_VOTER_wire)
  );
  defparam builder_array_muxed1_25_RED_VOTER.INIT = "0xFCC0";
  LUT4 builder_array_muxed1_26_RED_VOTER (
    .A(builder_array_muxed1_TMR_0[26]),
    .B(builder_array_muxed1_TMR_1[26]),
    .C(builder_array_muxed1_TMR_2[26]),
    .D(1'h0),
    .Z(builder_array_muxed1_26_RED_VOTER_wire)
  );
  defparam builder_array_muxed1_26_RED_VOTER.INIT = "0xFCC0";
  LUT4 builder_array_muxed1_27_RED_VOTER (
    .A(builder_array_muxed1_TMR_0[27]),
    .B(builder_array_muxed1_TMR_1[27]),
    .C(builder_array_muxed1_TMR_2[27]),
    .D(1'h0),
    .Z(builder_array_muxed1_27_RED_VOTER_wire)
  );
  defparam builder_array_muxed1_27_RED_VOTER.INIT = "0xFCC0";
  LUT4 builder_array_muxed1_28_RED_VOTER (
    .A(builder_array_muxed1_TMR_0[28]),
    .B(builder_array_muxed1_TMR_1[28]),
    .C(builder_array_muxed1_TMR_2[28]),
    .D(1'h0),
    .Z(builder_array_muxed1_28_RED_VOTER_wire)
  );
  defparam builder_array_muxed1_28_RED_VOTER.INIT = "0xFCC0";
  LUT4 builder_array_muxed1_29_RED_VOTER (
    .A(builder_array_muxed1_TMR_0[29]),
    .B(builder_array_muxed1_TMR_1[29]),
    .C(builder_array_muxed1_TMR_2[29]),
    .D(1'h0),
    .Z(builder_array_muxed1_29_RED_VOTER_wire)
  );
  defparam builder_array_muxed1_29_RED_VOTER.INIT = "0xFCC0";
  LUT4 builder_array_muxed1_2_RED_VOTER (
    .A(builder_array_muxed1_TMR_0[2]),
    .B(builder_array_muxed1_TMR_1[2]),
    .C(builder_array_muxed1_TMR_2[2]),
    .D(1'h0),
    .Z(builder_array_muxed1_2_RED_VOTER_wire)
  );
  defparam builder_array_muxed1_2_RED_VOTER.INIT = "0xFCC0";
  LUT4 builder_array_muxed1_30_RED_VOTER (
    .A(builder_array_muxed1_TMR_0[30]),
    .B(builder_array_muxed1_TMR_1[30]),
    .C(builder_array_muxed1_TMR_2[30]),
    .D(1'h0),
    .Z(builder_array_muxed1_30_RED_VOTER_wire)
  );
  defparam builder_array_muxed1_30_RED_VOTER.INIT = "0xFCC0";
  LUT4 builder_array_muxed1_31_RED_VOTER (
    .A(builder_array_muxed1_TMR_0[31]),
    .B(builder_array_muxed1_TMR_1[31]),
    .C(builder_array_muxed1_TMR_2[31]),
    .D(1'h0),
    .Z(builder_array_muxed1_31_RED_VOTER_wire)
  );
  defparam builder_array_muxed1_31_RED_VOTER.INIT = "0xFCC0";
  LUT4 builder_array_muxed1_3_RED_VOTER (
    .A(builder_array_muxed1_TMR_0[3]),
    .B(builder_array_muxed1_TMR_1[3]),
    .C(builder_array_muxed1_TMR_2[3]),
    .D(1'h0),
    .Z(builder_array_muxed1_3_RED_VOTER_wire)
  );
  defparam builder_array_muxed1_3_RED_VOTER.INIT = "0xFCC0";
  LUT4 builder_array_muxed1_4_RED_VOTER (
    .A(builder_array_muxed1_TMR_0[4]),
    .B(builder_array_muxed1_TMR_1[4]),
    .C(builder_array_muxed1_TMR_2[4]),
    .D(1'h0),
    .Z(builder_array_muxed1_4_RED_VOTER_wire)
  );
  defparam builder_array_muxed1_4_RED_VOTER.INIT = "0xFCC0";
  LUT4 builder_array_muxed1_5_RED_VOTER (
    .A(builder_array_muxed1_TMR_0[5]),
    .B(builder_array_muxed1_TMR_1[5]),
    .C(builder_array_muxed1_TMR_2[5]),
    .D(1'h0),
    .Z(builder_array_muxed1_5_RED_VOTER_wire)
  );
  defparam builder_array_muxed1_5_RED_VOTER.INIT = "0xFCC0";
  LUT4 builder_array_muxed1_6_RED_VOTER (
    .A(builder_array_muxed1_TMR_0[6]),
    .B(builder_array_muxed1_TMR_1[6]),
    .C(builder_array_muxed1_TMR_2[6]),
    .D(1'h0),
    .Z(builder_array_muxed1_6_RED_VOTER_wire)
  );
  defparam builder_array_muxed1_6_RED_VOTER.INIT = "0xFCC0";
  LUT4 builder_array_muxed1_7_RED_VOTER (
    .A(builder_array_muxed1_TMR_0[7]),
    .B(builder_array_muxed1_TMR_1[7]),
    .C(builder_array_muxed1_TMR_2[7]),
    .D(1'h0),
    .Z(builder_array_muxed1_7_RED_VOTER_wire)
  );
  defparam builder_array_muxed1_7_RED_VOTER.INIT = "0xFCC0";
  LUT4 builder_array_muxed1_8_RED_VOTER (
    .A(builder_array_muxed1_TMR_0[8]),
    .B(builder_array_muxed1_TMR_1[8]),
    .C(builder_array_muxed1_TMR_2[8]),
    .D(1'h0),
    .Z(builder_array_muxed1_8_RED_VOTER_wire)
  );
  defparam builder_array_muxed1_8_RED_VOTER.INIT = "0xFCC0";
  LUT4 builder_array_muxed1_9_RED_VOTER (
    .A(builder_array_muxed1_TMR_0[9]),
    .B(builder_array_muxed1_TMR_1[9]),
    .C(builder_array_muxed1_TMR_2[9]),
    .D(1'h0),
    .Z(builder_array_muxed1_9_RED_VOTER_wire)
  );
  defparam builder_array_muxed1_9_RED_VOTER.INIT = "0xFCC0";
  LUT4 builder_array_muxed2_i_0_RED_VOTER (
    .A(builder_array_muxed2_i_TMR_0[0]),
    .B(builder_array_muxed2_i_TMR_1[0]),
    .C(builder_array_muxed2_i_TMR_2[0]),
    .D(1'h0),
    .Z(builder_array_muxed2_i_0_RED_VOTER_wire)
  );
  defparam builder_array_muxed2_i_0_RED_VOTER.INIT = "0xFCC0";
  LUT4 builder_array_muxed2_i_1_RED_VOTER (
    .A(builder_array_muxed2_i_TMR_0[1]),
    .B(builder_array_muxed2_i_TMR_1[1]),
    .C(builder_array_muxed2_i_TMR_2[1]),
    .D(1'h0),
    .Z(builder_array_muxed2_i_1_RED_VOTER_wire)
  );
  defparam builder_array_muxed2_i_1_RED_VOTER.INIT = "0xFCC0";
  LUT4 builder_array_muxed2_i_2_RED_VOTER (
    .A(builder_array_muxed2_i_TMR_0[2]),
    .B(builder_array_muxed2_i_TMR_1[2]),
    .C(builder_array_muxed2_i_TMR_2[2]),
    .D(1'h0),
    .Z(builder_array_muxed2_i_2_RED_VOTER_wire)
  );
  defparam builder_array_muxed2_i_2_RED_VOTER.INIT = "0xFCC0";
  LUT4 builder_array_muxed2_i_3_RED_VOTER (
    .A(builder_array_muxed2_i_TMR_0[3]),
    .B(builder_array_muxed2_i_TMR_1[3]),
    .C(builder_array_muxed2_i_TMR_2[3]),
    .D(1'h0),
    .Z(builder_array_muxed2_i_3_RED_VOTER_wire)
  );
  defparam builder_array_muxed2_i_3_RED_VOTER.INIT = "0xFCC0";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51274.7-51277.2" *)
  INV builder_basesoc_rs232phyrx_state_RNISQ1C_TMR_0 (
    .A(builder_basesoc_rs232phyrx_state_TMR_0),
    .Z(builder_basesoc_rs232phyrx_state_i_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51274.7-51277.2" *)
  INV builder_basesoc_rs232phyrx_state_RNISQ1C_TMR_1 (
    .A(builder_basesoc_rs232phyrx_state_TMR_1),
    .Z(builder_basesoc_rs232phyrx_state_i_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51274.7-51277.2" *)
  INV builder_basesoc_rs232phyrx_state_RNISQ1C_TMR_2 (
    .A(builder_basesoc_rs232phyrx_state_TMR_2),
    .Z(builder_basesoc_rs232phyrx_state_i_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55485.11-55491.2" *)
  FD1P3IX builder_basesoc_rs232phyrx_state_reg_TMR_0 (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(N_110_TMR_0),
    .Q(builder_basesoc_rs232phyrx_state_TMR_0),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55485.11-55491.2" *)
  FD1P3IX builder_basesoc_rs232phyrx_state_reg_TMR_1 (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(N_110_TMR_1),
    .Q(builder_basesoc_rs232phyrx_state_TMR_1),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55485.11-55491.2" *)
  FD1P3IX builder_basesoc_rs232phyrx_state_reg_TMR_2 (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(N_110_TMR_2),
    .Q(builder_basesoc_rs232phyrx_state_TMR_2),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51269.7-51272.2" *)
  INV builder_basesoc_rs232phytx_state_RNIU8C3_TMR_0 (
    .A(builder_basesoc_rs232phytx_state_TMR_0),
    .Z(builder_basesoc_rs232phytx_state_i_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51269.7-51272.2" *)
  INV builder_basesoc_rs232phytx_state_RNIU8C3_TMR_1 (
    .A(builder_basesoc_rs232phytx_state_TMR_1),
    .Z(builder_basesoc_rs232phytx_state_i_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51269.7-51272.2" *)
  INV builder_basesoc_rs232phytx_state_RNIU8C3_TMR_2 (
    .A(builder_basesoc_rs232phytx_state_TMR_2),
    .Z(builder_basesoc_rs232phytx_state_i_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55478.11-55484.2" *)
  FD1P3IX builder_basesoc_rs232phytx_state_reg_TMR_0 (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(main_basesoc_tx_data_rs232phytx_next_value2_0_sqmuxa_TMR_0),
    .Q(builder_basesoc_rs232phytx_state_TMR_0),
    .SP(un1_main_basesoc_serial_tx_rs232phytx_next_value112_i_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55478.11-55484.2" *)
  FD1P3IX builder_basesoc_rs232phytx_state_reg_TMR_1 (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(main_basesoc_tx_data_rs232phytx_next_value2_0_sqmuxa_TMR_1),
    .Q(builder_basesoc_rs232phytx_state_TMR_1),
    .SP(un1_main_basesoc_serial_tx_rs232phytx_next_value112_i_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55478.11-55484.2" *)
  FD1P3IX builder_basesoc_rs232phytx_state_reg_TMR_2 (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(main_basesoc_tx_data_rs232phytx_next_value2_0_sqmuxa_TMR_2),
    .Q(builder_basesoc_rs232phytx_state_TMR_2),
    .SP(un1_main_basesoc_serial_tx_rs232phytx_next_value112_i_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55471.11-55477.2" *)
  FD1P3IX builder_basesoc_state_reg_TMR_0 (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_basesoc_next_state_1_sqmuxa_1_TMR_0),
    .Q(builder_basesoc_state_TMR_0),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55471.11-55477.2" *)
  FD1P3IX builder_basesoc_state_reg_TMR_1 (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_basesoc_next_state_1_sqmuxa_1_TMR_1),
    .Q(builder_basesoc_state_TMR_1),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55471.11-55477.2" *)
  FD1P3IX builder_basesoc_state_reg_TMR_2 (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_basesoc_next_state_1_sqmuxa_1_TMR_2),
    .Q(builder_basesoc_state_TMR_2),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55401.11-55407.2" *)
  FD1P3IX \builder_count[10]_TMR_0  (
    .CD(N_152_i_TMR_0),
    .CK(sys_clk),
    .D(builder_count_1_cry_9_0_S1_TMR_0),
    .Q(dsp_join_kb_25_TMR_0[10]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55401.11-55407.2" *)
  FD1P3IX \builder_count[10]_TMR_1  (
    .CD(N_152_i_TMR_1),
    .CK(sys_clk),
    .D(builder_count_1_cry_9_0_S1_TMR_1),
    .Q(dsp_join_kb_25_TMR_1[10]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55401.11-55407.2" *)
  FD1P3IX \builder_count[10]_TMR_2  (
    .CD(N_152_i_TMR_2),
    .CK(sys_clk),
    .D(builder_count_1_cry_9_0_S1_TMR_2),
    .Q(dsp_join_kb_25_TMR_2[10]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55408.11-55414.2" *)
  FD1P3IX \builder_count[11]_TMR_0  (
    .CD(N_152_i_TMR_0),
    .CK(sys_clk),
    .D(builder_count_1_cry_11_0_S0_TMR_0),
    .Q(dsp_join_kb_25_TMR_0[11]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55408.11-55414.2" *)
  FD1P3IX \builder_count[11]_TMR_1  (
    .CD(N_152_i_TMR_1),
    .CK(sys_clk),
    .D(builder_count_1_cry_11_0_S0_TMR_1),
    .Q(dsp_join_kb_25_TMR_1[11]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55408.11-55414.2" *)
  FD1P3IX \builder_count[11]_TMR_2  (
    .CD(N_152_i_TMR_2),
    .CK(sys_clk),
    .D(builder_count_1_cry_11_0_S0_TMR_2),
    .Q(dsp_join_kb_25_TMR_2[11]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55415.11-55421.2" *)
  FD1P3IX \builder_count[12]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_count_r_TMR_0[12]),
    .Q(dsp_join_kb_25_TMR_0[12]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55415.11-55421.2" *)
  FD1P3IX \builder_count[12]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_count_r_TMR_1[12]),
    .Q(dsp_join_kb_25_TMR_1[12]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55415.11-55421.2" *)
  FD1P3IX \builder_count[12]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_count_r_TMR_2[12]),
    .Q(dsp_join_kb_25_TMR_2[12]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55422.11-55428.2" *)
  FD1P3IX \builder_count[13]_TMR_0  (
    .CD(N_152_i_TMR_0),
    .CK(sys_clk),
    .D(builder_count_1_cry_13_0_S0_TMR_0),
    .Q(dsp_join_kb_25_TMR_0[13]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55422.11-55428.2" *)
  FD1P3IX \builder_count[13]_TMR_1  (
    .CD(N_152_i_TMR_1),
    .CK(sys_clk),
    .D(builder_count_1_cry_13_0_S0_TMR_1),
    .Q(dsp_join_kb_25_TMR_1[13]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55422.11-55428.2" *)
  FD1P3IX \builder_count[13]_TMR_2  (
    .CD(N_152_i_TMR_2),
    .CK(sys_clk),
    .D(builder_count_1_cry_13_0_S0_TMR_2),
    .Q(dsp_join_kb_25_TMR_2[13]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55429.11-55435.2" *)
  FD1P3JX \builder_count[14]_TMR_0  (
    .CK(sys_clk),
    .D(N_120_i_TMR_0),
    .PD(GND_0),
    .Q(dsp_join_kb_25_TMR_0[14]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55429.11-55435.2" *)
  FD1P3JX \builder_count[14]_TMR_1  (
    .CK(sys_clk),
    .D(N_120_i_TMR_1),
    .PD(GND_0),
    .Q(dsp_join_kb_25_TMR_1[14]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55429.11-55435.2" *)
  FD1P3JX \builder_count[14]_TMR_2  (
    .CK(sys_clk),
    .D(N_120_i_TMR_2),
    .PD(GND_0),
    .Q(dsp_join_kb_25_TMR_2[14]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55436.11-55442.2" *)
  FD1P3IX \builder_count[15]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_count_r_TMR_0[15]),
    .Q(dsp_join_kb_25_TMR_0[15]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55436.11-55442.2" *)
  FD1P3IX \builder_count[15]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_count_r_TMR_1[15]),
    .Q(dsp_join_kb_25_TMR_1[15]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55436.11-55442.2" *)
  FD1P3IX \builder_count[15]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_count_r_TMR_2[15]),
    .Q(dsp_join_kb_25_TMR_2[15]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55443.11-55449.2" *)
  FD1P3JX \builder_count[16]_TMR_0  (
    .CK(sys_clk),
    .D(N_121_i_TMR_0),
    .PD(GND_0),
    .Q(dsp_join_kb_25_TMR_0[16]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55443.11-55449.2" *)
  FD1P3JX \builder_count[16]_TMR_1  (
    .CK(sys_clk),
    .D(N_121_i_TMR_1),
    .PD(GND_0),
    .Q(dsp_join_kb_25_TMR_1[16]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55443.11-55449.2" *)
  FD1P3JX \builder_count[16]_TMR_2  (
    .CK(sys_clk),
    .D(N_121_i_TMR_2),
    .PD(GND_0),
    .Q(dsp_join_kb_25_TMR_2[16]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55450.11-55456.2" *)
  FD1P3JX \builder_count[17]_TMR_0  (
    .CK(sys_clk),
    .D(N_1218_i_TMR_0),
    .PD(GND_0),
    .Q(dsp_join_kb_25_TMR_0[17]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55450.11-55456.2" *)
  FD1P3JX \builder_count[17]_TMR_1  (
    .CK(sys_clk),
    .D(N_1218_i_TMR_1),
    .PD(GND_0),
    .Q(dsp_join_kb_25_TMR_1[17]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55450.11-55456.2" *)
  FD1P3JX \builder_count[17]_TMR_2  (
    .CK(sys_clk),
    .D(N_1218_i_TMR_2),
    .PD(GND_0),
    .Q(dsp_join_kb_25_TMR_2[17]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55457.11-55463.2" *)
  FD1P3JX \builder_count[18]_TMR_0  (
    .CK(sys_clk),
    .D(N_123_i_TMR_0),
    .PD(GND_0),
    .Q(dsp_join_kb_25_TMR_0[18]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55457.11-55463.2" *)
  FD1P3JX \builder_count[18]_TMR_1  (
    .CK(sys_clk),
    .D(N_123_i_TMR_1),
    .PD(GND_0),
    .Q(dsp_join_kb_25_TMR_1[18]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55457.11-55463.2" *)
  FD1P3JX \builder_count[18]_TMR_2  (
    .CK(sys_clk),
    .D(N_123_i_TMR_2),
    .PD(GND_0),
    .Q(dsp_join_kb_25_TMR_2[18]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55464.11-55470.2" *)
  FD1P3JX \builder_count[19]_TMR_0  (
    .CK(sys_clk),
    .D(N_124_i_TMR_0),
    .PD(GND_0),
    .Q(dsp_join_kb_25_TMR_0[19]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55464.11-55470.2" *)
  FD1P3JX \builder_count[19]_TMR_1  (
    .CK(sys_clk),
    .D(N_124_i_TMR_1),
    .PD(GND_0),
    .Q(dsp_join_kb_25_TMR_1[19]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55464.11-55470.2" *)
  FD1P3JX \builder_count[19]_TMR_2  (
    .CK(sys_clk),
    .D(N_124_i_TMR_2),
    .PD(GND_0),
    .Q(dsp_join_kb_25_TMR_2[19]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55373.11-55379.2" *)
  FD1P3JX \builder_count[6]_TMR_0  (
    .CK(sys_clk),
    .D(N_137_i_TMR_0),
    .PD(GND_0),
    .Q(dsp_join_kb_25_TMR_0[6]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55373.11-55379.2" *)
  FD1P3JX \builder_count[6]_TMR_1  (
    .CK(sys_clk),
    .D(N_137_i_TMR_1),
    .PD(GND_0),
    .Q(dsp_join_kb_25_TMR_1[6]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55373.11-55379.2" *)
  FD1P3JX \builder_count[6]_TMR_2  (
    .CK(sys_clk),
    .D(N_137_i_TMR_2),
    .PD(GND_0),
    .Q(dsp_join_kb_25_TMR_2[6]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55380.11-55386.2" *)
  FD1P3IX \builder_count[7]_TMR_0  (
    .CD(N_152_i_TMR_0),
    .CK(sys_clk),
    .D(builder_count_1_cry_7_0_S0_TMR_0),
    .Q(dsp_join_kb_25_TMR_0[7]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55380.11-55386.2" *)
  FD1P3IX \builder_count[7]_TMR_1  (
    .CD(N_152_i_TMR_1),
    .CK(sys_clk),
    .D(builder_count_1_cry_7_0_S0_TMR_1),
    .Q(dsp_join_kb_25_TMR_1[7]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55380.11-55386.2" *)
  FD1P3IX \builder_count[7]_TMR_2  (
    .CD(N_152_i_TMR_2),
    .CK(sys_clk),
    .D(builder_count_1_cry_7_0_S0_TMR_2),
    .Q(dsp_join_kb_25_TMR_2[7]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55387.11-55393.2" *)
  FD1P3IX \builder_count[8]_TMR_0  (
    .CD(N_152_i_TMR_0),
    .CK(sys_clk),
    .D(builder_count_1_cry_7_0_S1_TMR_0),
    .Q(dsp_join_kb_25_TMR_0[8]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55387.11-55393.2" *)
  FD1P3IX \builder_count[8]_TMR_1  (
    .CD(N_152_i_TMR_1),
    .CK(sys_clk),
    .D(builder_count_1_cry_7_0_S1_TMR_1),
    .Q(dsp_join_kb_25_TMR_1[8]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55387.11-55393.2" *)
  FD1P3IX \builder_count[8]_TMR_2  (
    .CD(N_152_i_TMR_2),
    .CK(sys_clk),
    .D(builder_count_1_cry_7_0_S1_TMR_2),
    .Q(dsp_join_kb_25_TMR_2[8]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55394.11-55400.2" *)
  FD1P3JX \builder_count[9]_TMR_0  (
    .CK(sys_clk),
    .D(N_1219_i_TMR_0),
    .PD(GND_0),
    .Q(dsp_join_kb_25_TMR_0[9]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55394.11-55400.2" *)
  FD1P3JX \builder_count[9]_TMR_1  (
    .CK(sys_clk),
    .D(N_1219_i_TMR_1),
    .PD(GND_0),
    .Q(dsp_join_kb_25_TMR_1[9]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55394.11-55400.2" *)
  FD1P3JX \builder_count[9]_TMR_2  (
    .CK(sys_clk),
    .D(N_1219_i_TMR_2),
    .PD(GND_0),
    .Q(dsp_join_kb_25_TMR_2[9]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55345.11-55351.2" *)
  FD1P3IX \builder_count_0_mod[0]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_count_0_mod_RNO_TMR_0[0]),
    .Q(builder_count_1_TMR_0),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55345.11-55351.2" *)
  FD1P3IX \builder_count_0_mod[0]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_count_0_mod_RNO_TMR_1[0]),
    .Q(builder_count_1_TMR_1),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55345.11-55351.2" *)
  FD1P3IX \builder_count_0_mod[0]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_count_0_mod_RNO_TMR_2[0]),
    .Q(builder_count_1_TMR_2),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55352.11-55358.2" *)
  FD1P3IX \builder_count_0_mod[1]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_count_0_mod_RNO_TMR_0[1]),
    .Q(dsp_join_kb_25_TMR_0[1]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55352.11-55358.2" *)
  FD1P3IX \builder_count_0_mod[1]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_count_0_mod_RNO_TMR_1[1]),
    .Q(dsp_join_kb_25_TMR_1[1]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55352.11-55358.2" *)
  FD1P3IX \builder_count_0_mod[1]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_count_0_mod_RNO_TMR_2[1]),
    .Q(dsp_join_kb_25_TMR_2[1]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55359.11-55365.2" *)
  FD1P3IX \builder_count_0_mod[3]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_count_0_mod_RNO_TMR_0[3]),
    .Q(dsp_join_kb_25_TMR_0[3]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55359.11-55365.2" *)
  FD1P3IX \builder_count_0_mod[3]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_count_0_mod_RNO_TMR_1[3]),
    .Q(dsp_join_kb_25_TMR_1[3]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55359.11-55365.2" *)
  FD1P3IX \builder_count_0_mod[3]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_count_0_mod_RNO_TMR_2[3]),
    .Q(dsp_join_kb_25_TMR_2[3]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55366.11-55372.2" *)
  FD1P3IX \builder_count_0_mod[5]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_count_0_mod_RNO_TMR_0[5]),
    .Q(dsp_join_kb_25_TMR_0[5]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55366.11-55372.2" *)
  FD1P3IX \builder_count_0_mod[5]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_count_0_mod_RNO_TMR_1[5]),
    .Q(dsp_join_kb_25_TMR_1[5]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55366.11-55372.2" *)
  FD1P3IX \builder_count_0_mod[5]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_count_0_mod_RNO_TMR_2[5]),
    .Q(dsp_join_kb_25_TMR_2[5]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51326.8-51332.2" *)
  LUT4 \builder_count_0_mod_RNO_cZ[0]_TMR_0  (
    .A(builder_count_1_TMR_0),
    .B(builder_wait_TMR_0),
    .C(sys_rst_TMR_0),
    .D(GND_0),
    .Z(builder_count_0_mod_RNO_TMR_0[0])
  );
  defparam \builder_count_0_mod_RNO_cZ[0]_TMR_0 .INIT = "0x0404";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51326.8-51332.2" *)
  LUT4 \builder_count_0_mod_RNO_cZ[0]_TMR_1  (
    .A(builder_count_1_TMR_1),
    .B(builder_wait_TMR_1),
    .C(sys_rst_TMR_1),
    .D(GND_0),
    .Z(builder_count_0_mod_RNO_TMR_1[0])
  );
  defparam \builder_count_0_mod_RNO_cZ[0]_TMR_1 .INIT = "0x0404";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51326.8-51332.2" *)
  LUT4 \builder_count_0_mod_RNO_cZ[0]_TMR_2  (
    .A(builder_count_1_TMR_2),
    .B(builder_wait_TMR_2),
    .C(sys_rst_TMR_2),
    .D(GND_0),
    .Z(builder_count_0_mod_RNO_TMR_2[0])
  );
  defparam \builder_count_0_mod_RNO_cZ[0]_TMR_2 .INIT = "0x0404";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51317.8-51323.2" *)
  LUT4 \builder_count_0_mod_RNO_cZ[1]_TMR_0  (
    .A(builder_count_1_cry_1_0_S0_TMR_0),
    .B(builder_wait_TMR_0),
    .C(sys_rst_TMR_0),
    .D(GND_0),
    .Z(builder_count_0_mod_RNO_TMR_0[1])
  );
  defparam \builder_count_0_mod_RNO_cZ[1]_TMR_0 .INIT = "0x0808";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51317.8-51323.2" *)
  LUT4 \builder_count_0_mod_RNO_cZ[1]_TMR_1  (
    .A(builder_count_1_cry_1_0_S0_TMR_1),
    .B(builder_wait_TMR_1),
    .C(sys_rst_TMR_1),
    .D(GND_0),
    .Z(builder_count_0_mod_RNO_TMR_1[1])
  );
  defparam \builder_count_0_mod_RNO_cZ[1]_TMR_1 .INIT = "0x0808";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51317.8-51323.2" *)
  LUT4 \builder_count_0_mod_RNO_cZ[1]_TMR_2  (
    .A(builder_count_1_cry_1_0_S0_TMR_2),
    .B(builder_wait_TMR_2),
    .C(sys_rst_TMR_2),
    .D(GND_0),
    .Z(builder_count_0_mod_RNO_TMR_2[1])
  );
  defparam \builder_count_0_mod_RNO_cZ[1]_TMR_2 .INIT = "0x0808";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51308.8-51314.2" *)
  LUT4 \builder_count_0_mod_RNO_cZ[3]_TMR_0  (
    .A(N_698_TMR_0),
    .B(builder_wait_TMR_0),
    .C(sys_rst_TMR_0),
    .D(GND_0),
    .Z(builder_count_0_mod_RNO_TMR_0[3])
  );
  defparam \builder_count_0_mod_RNO_cZ[3]_TMR_0 .INIT = "0x0808";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51308.8-51314.2" *)
  LUT4 \builder_count_0_mod_RNO_cZ[3]_TMR_1  (
    .A(N_698_TMR_1),
    .B(builder_wait_TMR_1),
    .C(sys_rst_TMR_1),
    .D(GND_0),
    .Z(builder_count_0_mod_RNO_TMR_1[3])
  );
  defparam \builder_count_0_mod_RNO_cZ[3]_TMR_1 .INIT = "0x0808";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51308.8-51314.2" *)
  LUT4 \builder_count_0_mod_RNO_cZ[3]_TMR_2  (
    .A(N_698_TMR_2),
    .B(builder_wait_TMR_2),
    .C(sys_rst_TMR_2),
    .D(GND_0),
    .Z(builder_count_0_mod_RNO_TMR_2[3])
  );
  defparam \builder_count_0_mod_RNO_cZ[3]_TMR_2 .INIT = "0x0808";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51299.8-51305.2" *)
  LUT4 \builder_count_0_mod_RNO_cZ[5]_TMR_0  (
    .A(builder_count_1_cry_5_0_S0_TMR_0),
    .B(builder_wait_TMR_0),
    .C(sys_rst_TMR_0),
    .D(GND_0),
    .Z(builder_count_0_mod_RNO_TMR_0[5])
  );
  defparam \builder_count_0_mod_RNO_cZ[5]_TMR_0 .INIT = "0x0808";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51299.8-51305.2" *)
  LUT4 \builder_count_0_mod_RNO_cZ[5]_TMR_1  (
    .A(builder_count_1_cry_5_0_S0_TMR_1),
    .B(builder_wait_TMR_1),
    .C(sys_rst_TMR_1),
    .D(GND_0),
    .Z(builder_count_0_mod_RNO_TMR_1[5])
  );
  defparam \builder_count_0_mod_RNO_cZ[5]_TMR_1 .INIT = "0x0808";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51299.8-51305.2" *)
  LUT4 \builder_count_0_mod_RNO_cZ[5]_TMR_2  (
    .A(builder_count_1_cry_5_0_S0_TMR_2),
    .B(builder_wait_TMR_2),
    .C(sys_rst_TMR_2),
    .D(GND_0),
    .Z(builder_count_0_mod_RNO_TMR_2[5])
  );
  defparam \builder_count_0_mod_RNO_cZ[5]_TMR_2 .INIT = "0x0808";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57714.8-57727.2" *)
  CCU2 builder_count_1_cry_0_0_TMR_0 (
    .A0(VCC_TMR_0),
    .A1(builder_count_1_TMR_0),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(GND_0),
    .COUT(builder_count_1_cry_0_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(builder_count_1_cry_0_0_S0_TMR_0),
    .S1(builder_count_1_cry_0_0_S1_TMR_0)
  );
  defparam builder_count_1_cry_0_0_TMR_0.INIT0 = "5033";
  defparam builder_count_1_cry_0_0_TMR_0.INIT1 = "50AA";
  defparam builder_count_1_cry_0_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57714.8-57727.2" *)
  CCU2 builder_count_1_cry_0_0_TMR_1 (
    .A0(VCC_TMR_1),
    .A1(builder_count_1_TMR_1),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(GND_0),
    .COUT(builder_count_1_cry_0_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(builder_count_1_cry_0_0_S0_TMR_1),
    .S1(builder_count_1_cry_0_0_S1_TMR_1)
  );
  defparam builder_count_1_cry_0_0_TMR_1.INIT0 = "5033";
  defparam builder_count_1_cry_0_0_TMR_1.INIT1 = "50AA";
  defparam builder_count_1_cry_0_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57714.8-57727.2" *)
  CCU2 builder_count_1_cry_0_0_TMR_2 (
    .A0(VCC_TMR_2),
    .A1(builder_count_1_TMR_2),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(GND_0),
    .COUT(builder_count_1_cry_0_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(builder_count_1_cry_0_0_S0_TMR_2),
    .S1(builder_count_1_cry_0_0_S1_TMR_2)
  );
  defparam builder_count_1_cry_0_0_TMR_2.INIT0 = "5033";
  defparam builder_count_1_cry_0_0_TMR_2.INIT1 = "50AA";
  defparam builder_count_1_cry_0_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57607.8-57620.2" *)
  CCU2 builder_count_1_cry_11_0_TMR_0 (
    .A0(dsp_join_kb_25_TMR_0[11]),
    .A1(dsp_join_kb_25_TMR_0[12]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(builder_count_1_cry_10_TMR_0),
    .COUT(builder_count_1_cry_12_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(builder_count_1_cry_11_0_S0_TMR_0),
    .S1(builder_count_1_cry_11_0_S1_TMR_0)
  );
  defparam builder_count_1_cry_11_0_TMR_0.INIT0 = "50AA";
  defparam builder_count_1_cry_11_0_TMR_0.INIT1 = "50AA";
  defparam builder_count_1_cry_11_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57607.8-57620.2" *)
  CCU2 builder_count_1_cry_11_0_TMR_1 (
    .A0(dsp_join_kb_25_TMR_1[11]),
    .A1(dsp_join_kb_25_TMR_1[12]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(builder_count_1_cry_10_TMR_1),
    .COUT(builder_count_1_cry_12_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(builder_count_1_cry_11_0_S0_TMR_1),
    .S1(builder_count_1_cry_11_0_S1_TMR_1)
  );
  defparam builder_count_1_cry_11_0_TMR_1.INIT0 = "50AA";
  defparam builder_count_1_cry_11_0_TMR_1.INIT1 = "50AA";
  defparam builder_count_1_cry_11_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57607.8-57620.2" *)
  CCU2 builder_count_1_cry_11_0_TMR_2 (
    .A0(dsp_join_kb_25_TMR_2[11]),
    .A1(dsp_join_kb_25_TMR_2[12]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(builder_count_1_cry_10_TMR_2),
    .COUT(builder_count_1_cry_12_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(builder_count_1_cry_11_0_S0_TMR_2),
    .S1(builder_count_1_cry_11_0_S1_TMR_2)
  );
  defparam builder_count_1_cry_11_0_TMR_2.INIT0 = "50AA";
  defparam builder_count_1_cry_11_0_TMR_2.INIT1 = "50AA";
  defparam builder_count_1_cry_11_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57589.8-57602.2" *)
  CCU2 builder_count_1_cry_13_0_TMR_0 (
    .A0(dsp_join_kb_25_TMR_0[13]),
    .A1(dsp_join_kb_25_TMR_0[14]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(builder_count_1_cry_12_TMR_0),
    .COUT(builder_count_1_cry_14_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(builder_count_1_cry_13_0_S0_TMR_0),
    .S1(builder_count_1_2_TMR_0[14])
  );
  defparam builder_count_1_cry_13_0_TMR_0.INIT0 = "50AA";
  defparam builder_count_1_cry_13_0_TMR_0.INIT1 = "50AA";
  defparam builder_count_1_cry_13_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57589.8-57602.2" *)
  CCU2 builder_count_1_cry_13_0_TMR_1 (
    .A0(dsp_join_kb_25_TMR_1[13]),
    .A1(dsp_join_kb_25_TMR_1[14]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(builder_count_1_cry_12_TMR_1),
    .COUT(builder_count_1_cry_14_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(builder_count_1_cry_13_0_S0_TMR_1),
    .S1(builder_count_1_2_TMR_1[14])
  );
  defparam builder_count_1_cry_13_0_TMR_1.INIT0 = "50AA";
  defparam builder_count_1_cry_13_0_TMR_1.INIT1 = "50AA";
  defparam builder_count_1_cry_13_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57589.8-57602.2" *)
  CCU2 builder_count_1_cry_13_0_TMR_2 (
    .A0(dsp_join_kb_25_TMR_2[13]),
    .A1(dsp_join_kb_25_TMR_2[14]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(builder_count_1_cry_12_TMR_2),
    .COUT(builder_count_1_cry_14_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(builder_count_1_cry_13_0_S0_TMR_2),
    .S1(builder_count_1_2_TMR_2[14])
  );
  defparam builder_count_1_cry_13_0_TMR_2.INIT0 = "50AA";
  defparam builder_count_1_cry_13_0_TMR_2.INIT1 = "50AA";
  defparam builder_count_1_cry_13_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57571.8-57584.2" *)
  CCU2 builder_count_1_cry_15_0_TMR_0 (
    .A0(dsp_join_kb_25_TMR_0[15]),
    .A1(dsp_join_kb_25_TMR_0[16]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(builder_count_1_cry_14_TMR_0),
    .COUT(builder_count_1_cry_16_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(builder_count_1_cry_15_0_S0_TMR_0),
    .S1(builder_count_1_2_TMR_0[16])
  );
  defparam builder_count_1_cry_15_0_TMR_0.INIT0 = "50AA";
  defparam builder_count_1_cry_15_0_TMR_0.INIT1 = "50AA";
  defparam builder_count_1_cry_15_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57571.8-57584.2" *)
  CCU2 builder_count_1_cry_15_0_TMR_1 (
    .A0(dsp_join_kb_25_TMR_1[15]),
    .A1(dsp_join_kb_25_TMR_1[16]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(builder_count_1_cry_14_TMR_1),
    .COUT(builder_count_1_cry_16_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(builder_count_1_cry_15_0_S0_TMR_1),
    .S1(builder_count_1_2_TMR_1[16])
  );
  defparam builder_count_1_cry_15_0_TMR_1.INIT0 = "50AA";
  defparam builder_count_1_cry_15_0_TMR_1.INIT1 = "50AA";
  defparam builder_count_1_cry_15_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57571.8-57584.2" *)
  CCU2 builder_count_1_cry_15_0_TMR_2 (
    .A0(dsp_join_kb_25_TMR_2[15]),
    .A1(dsp_join_kb_25_TMR_2[16]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(builder_count_1_cry_14_TMR_2),
    .COUT(builder_count_1_cry_16_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(builder_count_1_cry_15_0_S0_TMR_2),
    .S1(builder_count_1_2_TMR_2[16])
  );
  defparam builder_count_1_cry_15_0_TMR_2.INIT0 = "50AA";
  defparam builder_count_1_cry_15_0_TMR_2.INIT1 = "50AA";
  defparam builder_count_1_cry_15_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57553.8-57566.2" *)
  CCU2 builder_count_1_cry_17_0_TMR_0 (
    .A0(dsp_join_kb_25_TMR_0[17]),
    .A1(dsp_join_kb_25_TMR_0[18]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(builder_count_1_cry_16_TMR_0),
    .COUT(builder_count_1_cry_18_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(builder_count_1_2_TMR_0[17]),
    .S1(builder_count_1_2_TMR_0[18])
  );
  defparam builder_count_1_cry_17_0_TMR_0.INIT0 = "50AA";
  defparam builder_count_1_cry_17_0_TMR_0.INIT1 = "50FF";
  defparam builder_count_1_cry_17_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57553.8-57566.2" *)
  CCU2 builder_count_1_cry_17_0_TMR_1 (
    .A0(dsp_join_kb_25_TMR_1[17]),
    .A1(dsp_join_kb_25_TMR_1[18]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(builder_count_1_cry_16_TMR_1),
    .COUT(builder_count_1_cry_18_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(builder_count_1_2_TMR_1[17]),
    .S1(builder_count_1_2_TMR_1[18])
  );
  defparam builder_count_1_cry_17_0_TMR_1.INIT0 = "50AA";
  defparam builder_count_1_cry_17_0_TMR_1.INIT1 = "50FF";
  defparam builder_count_1_cry_17_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57553.8-57566.2" *)
  CCU2 builder_count_1_cry_17_0_TMR_2 (
    .A0(dsp_join_kb_25_TMR_2[17]),
    .A1(dsp_join_kb_25_TMR_2[18]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(builder_count_1_cry_16_TMR_2),
    .COUT(builder_count_1_cry_18_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(builder_count_1_2_TMR_2[17]),
    .S1(builder_count_1_2_TMR_2[18])
  );
  defparam builder_count_1_cry_17_0_TMR_2.INIT0 = "50AA";
  defparam builder_count_1_cry_17_0_TMR_2.INIT1 = "50FF";
  defparam builder_count_1_cry_17_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57697.8-57710.2" *)
  CCU2 builder_count_1_cry_1_0_TMR_0 (
    .A0(dsp_join_kb_25_TMR_0[1]),
    .A1(dsp_join_kb_25_TMR_0[2]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(builder_count_1_cry_0_TMR_0),
    .COUT(builder_count_1_cry_2_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(builder_count_1_cry_1_0_S0_TMR_0),
    .S1(N_697_TMR_0)
  );
  defparam builder_count_1_cry_1_0_TMR_0.INIT0 = "50AA";
  defparam builder_count_1_cry_1_0_TMR_0.INIT1 = "50AA";
  defparam builder_count_1_cry_1_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57697.8-57710.2" *)
  CCU2 builder_count_1_cry_1_0_TMR_1 (
    .A0(dsp_join_kb_25_TMR_1[1]),
    .A1(dsp_join_kb_25_TMR_1[2]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(builder_count_1_cry_0_TMR_1),
    .COUT(builder_count_1_cry_2_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(builder_count_1_cry_1_0_S0_TMR_1),
    .S1(N_697_TMR_1)
  );
  defparam builder_count_1_cry_1_0_TMR_1.INIT0 = "50AA";
  defparam builder_count_1_cry_1_0_TMR_1.INIT1 = "50AA";
  defparam builder_count_1_cry_1_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57697.8-57710.2" *)
  CCU2 builder_count_1_cry_1_0_TMR_2 (
    .A0(dsp_join_kb_25_TMR_2[1]),
    .A1(dsp_join_kb_25_TMR_2[2]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(builder_count_1_cry_0_TMR_2),
    .COUT(builder_count_1_cry_2_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(builder_count_1_cry_1_0_S0_TMR_2),
    .S1(N_697_TMR_2)
  );
  defparam builder_count_1_cry_1_0_TMR_2.INIT0 = "50AA";
  defparam builder_count_1_cry_1_0_TMR_2.INIT1 = "50AA";
  defparam builder_count_1_cry_1_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57679.8-57692.2" *)
  CCU2 builder_count_1_cry_3_0_TMR_0 (
    .A0(dsp_join_kb_25_TMR_0[3]),
    .A1(dsp_join_kb_25_TMR_0[4]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(builder_count_1_cry_2_TMR_0),
    .COUT(builder_count_1_cry_4_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(N_698_TMR_0),
    .S1(N_699_TMR_0)
  );
  defparam builder_count_1_cry_3_0_TMR_0.INIT0 = "50AA";
  defparam builder_count_1_cry_3_0_TMR_0.INIT1 = "50AA";
  defparam builder_count_1_cry_3_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57679.8-57692.2" *)
  CCU2 builder_count_1_cry_3_0_TMR_1 (
    .A0(dsp_join_kb_25_TMR_1[3]),
    .A1(dsp_join_kb_25_TMR_1[4]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(builder_count_1_cry_2_TMR_1),
    .COUT(builder_count_1_cry_4_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(N_698_TMR_1),
    .S1(N_699_TMR_1)
  );
  defparam builder_count_1_cry_3_0_TMR_1.INIT0 = "50AA";
  defparam builder_count_1_cry_3_0_TMR_1.INIT1 = "50AA";
  defparam builder_count_1_cry_3_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57679.8-57692.2" *)
  CCU2 builder_count_1_cry_3_0_TMR_2 (
    .A0(dsp_join_kb_25_TMR_2[3]),
    .A1(dsp_join_kb_25_TMR_2[4]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(builder_count_1_cry_2_TMR_2),
    .COUT(builder_count_1_cry_4_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(N_698_TMR_2),
    .S1(N_699_TMR_2)
  );
  defparam builder_count_1_cry_3_0_TMR_2.INIT0 = "50AA";
  defparam builder_count_1_cry_3_0_TMR_2.INIT1 = "50AA";
  defparam builder_count_1_cry_3_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57661.8-57674.2" *)
  CCU2 builder_count_1_cry_5_0_TMR_0 (
    .A0(dsp_join_kb_25_TMR_0[5]),
    .A1(dsp_join_kb_25_TMR_0[6]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(builder_count_1_cry_4_TMR_0),
    .COUT(builder_count_1_cry_6_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(builder_count_1_cry_5_0_S0_TMR_0),
    .S1(builder_count_1_2_TMR_0[6])
  );
  defparam builder_count_1_cry_5_0_TMR_0.INIT0 = "50AA";
  defparam builder_count_1_cry_5_0_TMR_0.INIT1 = "50AA";
  defparam builder_count_1_cry_5_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57661.8-57674.2" *)
  CCU2 builder_count_1_cry_5_0_TMR_1 (
    .A0(dsp_join_kb_25_TMR_1[5]),
    .A1(dsp_join_kb_25_TMR_1[6]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(builder_count_1_cry_4_TMR_1),
    .COUT(builder_count_1_cry_6_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(builder_count_1_cry_5_0_S0_TMR_1),
    .S1(builder_count_1_2_TMR_1[6])
  );
  defparam builder_count_1_cry_5_0_TMR_1.INIT0 = "50AA";
  defparam builder_count_1_cry_5_0_TMR_1.INIT1 = "50AA";
  defparam builder_count_1_cry_5_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57661.8-57674.2" *)
  CCU2 builder_count_1_cry_5_0_TMR_2 (
    .A0(dsp_join_kb_25_TMR_2[5]),
    .A1(dsp_join_kb_25_TMR_2[6]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(builder_count_1_cry_4_TMR_2),
    .COUT(builder_count_1_cry_6_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(builder_count_1_cry_5_0_S0_TMR_2),
    .S1(builder_count_1_2_TMR_2[6])
  );
  defparam builder_count_1_cry_5_0_TMR_2.INIT0 = "50AA";
  defparam builder_count_1_cry_5_0_TMR_2.INIT1 = "50AA";
  defparam builder_count_1_cry_5_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57643.8-57656.2" *)
  CCU2 builder_count_1_cry_7_0_TMR_0 (
    .A0(dsp_join_kb_25_TMR_0[7]),
    .A1(dsp_join_kb_25_TMR_0[8]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(builder_count_1_cry_6_TMR_0),
    .COUT(builder_count_1_cry_8_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(builder_count_1_cry_7_0_S0_TMR_0),
    .S1(builder_count_1_cry_7_0_S1_TMR_0)
  );
  defparam builder_count_1_cry_7_0_TMR_0.INIT0 = "50AA";
  defparam builder_count_1_cry_7_0_TMR_0.INIT1 = "50AA";
  defparam builder_count_1_cry_7_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57643.8-57656.2" *)
  CCU2 builder_count_1_cry_7_0_TMR_1 (
    .A0(dsp_join_kb_25_TMR_1[7]),
    .A1(dsp_join_kb_25_TMR_1[8]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(builder_count_1_cry_6_TMR_1),
    .COUT(builder_count_1_cry_8_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(builder_count_1_cry_7_0_S0_TMR_1),
    .S1(builder_count_1_cry_7_0_S1_TMR_1)
  );
  defparam builder_count_1_cry_7_0_TMR_1.INIT0 = "50AA";
  defparam builder_count_1_cry_7_0_TMR_1.INIT1 = "50AA";
  defparam builder_count_1_cry_7_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57643.8-57656.2" *)
  CCU2 builder_count_1_cry_7_0_TMR_2 (
    .A0(dsp_join_kb_25_TMR_2[7]),
    .A1(dsp_join_kb_25_TMR_2[8]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(builder_count_1_cry_6_TMR_2),
    .COUT(builder_count_1_cry_8_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(builder_count_1_cry_7_0_S0_TMR_2),
    .S1(builder_count_1_cry_7_0_S1_TMR_2)
  );
  defparam builder_count_1_cry_7_0_TMR_2.INIT0 = "50AA";
  defparam builder_count_1_cry_7_0_TMR_2.INIT1 = "50AA";
  defparam builder_count_1_cry_7_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57625.8-57638.2" *)
  CCU2 builder_count_1_cry_9_0_TMR_0 (
    .A0(dsp_join_kb_25_TMR_0[9]),
    .A1(dsp_join_kb_25_TMR_0[10]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(builder_count_1_cry_8_TMR_0),
    .COUT(builder_count_1_cry_10_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(builder_count_1_2_TMR_0[9]),
    .S1(builder_count_1_cry_9_0_S1_TMR_0)
  );
  defparam builder_count_1_cry_9_0_TMR_0.INIT0 = "50AA";
  defparam builder_count_1_cry_9_0_TMR_0.INIT1 = "50AA";
  defparam builder_count_1_cry_9_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57625.8-57638.2" *)
  CCU2 builder_count_1_cry_9_0_TMR_1 (
    .A0(dsp_join_kb_25_TMR_1[9]),
    .A1(dsp_join_kb_25_TMR_1[10]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(builder_count_1_cry_8_TMR_1),
    .COUT(builder_count_1_cry_10_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(builder_count_1_2_TMR_1[9]),
    .S1(builder_count_1_cry_9_0_S1_TMR_1)
  );
  defparam builder_count_1_cry_9_0_TMR_1.INIT0 = "50AA";
  defparam builder_count_1_cry_9_0_TMR_1.INIT1 = "50AA";
  defparam builder_count_1_cry_9_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57625.8-57638.2" *)
  CCU2 builder_count_1_cry_9_0_TMR_2 (
    .A0(dsp_join_kb_25_TMR_2[9]),
    .A1(dsp_join_kb_25_TMR_2[10]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(builder_count_1_cry_8_TMR_2),
    .COUT(builder_count_1_cry_10_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(builder_count_1_2_TMR_2[9]),
    .S1(builder_count_1_cry_9_0_S1_TMR_2)
  );
  defparam builder_count_1_cry_9_0_TMR_2.INIT0 = "50AA";
  defparam builder_count_1_cry_9_0_TMR_2.INIT1 = "50AA";
  defparam builder_count_1_cry_9_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51289.7-51292.2" *)
  INV builder_count_1_s_19_0_RNO_TMR_0 (
    .A(dsp_join_kb_25_TMR_0[19]),
    .Z(dsp_join_kb_25_i_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51289.7-51292.2" *)
  INV builder_count_1_s_19_0_RNO_TMR_1 (
    .A(dsp_join_kb_25_TMR_1[19]),
    .Z(dsp_join_kb_25_i_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51289.7-51292.2" *)
  INV builder_count_1_s_19_0_RNO_TMR_2 (
    .A(dsp_join_kb_25_TMR_2[19]),
    .Z(dsp_join_kb_25_i_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57535.8-57548.2" *)
  CCU2 builder_count_1_s_19_0_TMR_0 (
    .A0(dsp_join_kb_25_i_TMR_0),
    .A1(VCC_TMR_0),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(builder_count_1_cry_18_TMR_0),
    .COUT(builder_count_1_s_19_0_COUT_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(builder_count_1_2_TMR_0[19]),
    .S1(builder_count_1_s_19_0_S1_TMR_0)
  );
  defparam builder_count_1_s_19_0_TMR_0.INIT0 = "A033";
  defparam builder_count_1_s_19_0_TMR_0.INIT1 = "5033";
  defparam builder_count_1_s_19_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57535.8-57548.2" *)
  CCU2 builder_count_1_s_19_0_TMR_1 (
    .A0(dsp_join_kb_25_i_TMR_1),
    .A1(VCC_TMR_1),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(builder_count_1_cry_18_TMR_1),
    .COUT(builder_count_1_s_19_0_COUT_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(builder_count_1_2_TMR_1[19]),
    .S1(builder_count_1_s_19_0_S1_TMR_1)
  );
  defparam builder_count_1_s_19_0_TMR_1.INIT0 = "A033";
  defparam builder_count_1_s_19_0_TMR_1.INIT1 = "5033";
  defparam builder_count_1_s_19_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57535.8-57548.2" *)
  CCU2 builder_count_1_s_19_0_TMR_2 (
    .A0(dsp_join_kb_25_i_TMR_2),
    .A1(VCC_TMR_2),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(builder_count_1_cry_18_TMR_2),
    .COUT(builder_count_1_s_19_0_COUT_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(builder_count_1_2_TMR_2[19]),
    .S1(builder_count_1_s_19_0_S1_TMR_2)
  );
  defparam builder_count_1_s_19_0_TMR_2.INIT0 = "A033";
  defparam builder_count_1_s_19_0_TMR_2.INIT1 = "5033";
  defparam builder_count_1_s_19_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55331.11-55337.2" *)
  FD1P3IX \builder_count_mod[2]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_count_mod_RNO_TMR_0[2]),
    .Q(dsp_join_kb_25_TMR_0[2]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55331.11-55337.2" *)
  FD1P3IX \builder_count_mod[2]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_count_mod_RNO_TMR_1[2]),
    .Q(dsp_join_kb_25_TMR_1[2]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55331.11-55337.2" *)
  FD1P3IX \builder_count_mod[2]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_count_mod_RNO_TMR_2[2]),
    .Q(dsp_join_kb_25_TMR_2[2]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55338.11-55344.2" *)
  FD1P3IX \builder_count_mod[4]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_count_mod_RNO_TMR_0[4]),
    .Q(dsp_join_kb_25_TMR_0[4]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55338.11-55344.2" *)
  FD1P3IX \builder_count_mod[4]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_count_mod_RNO_TMR_1[4]),
    .Q(dsp_join_kb_25_TMR_1[4]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55338.11-55344.2" *)
  FD1P3IX \builder_count_mod[4]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_count_mod_RNO_TMR_2[4]),
    .Q(dsp_join_kb_25_TMR_2[4]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51344.8-51350.2" *)
  LUT4 \builder_count_mod_RNO_cZ[2]_TMR_0  (
    .A(N_697_TMR_0),
    .B(builder_wait_TMR_0),
    .C(sys_rst_TMR_0),
    .D(GND_0),
    .Z(builder_count_mod_RNO_TMR_0[2])
  );
  defparam \builder_count_mod_RNO_cZ[2]_TMR_0 .INIT = "0x0808";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51344.8-51350.2" *)
  LUT4 \builder_count_mod_RNO_cZ[2]_TMR_1  (
    .A(N_697_TMR_1),
    .B(builder_wait_TMR_1),
    .C(sys_rst_TMR_1),
    .D(GND_0),
    .Z(builder_count_mod_RNO_TMR_1[2])
  );
  defparam \builder_count_mod_RNO_cZ[2]_TMR_1 .INIT = "0x0808";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51344.8-51350.2" *)
  LUT4 \builder_count_mod_RNO_cZ[2]_TMR_2  (
    .A(N_697_TMR_2),
    .B(builder_wait_TMR_2),
    .C(sys_rst_TMR_2),
    .D(GND_0),
    .Z(builder_count_mod_RNO_TMR_2[2])
  );
  defparam \builder_count_mod_RNO_cZ[2]_TMR_2 .INIT = "0x0808";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51335.8-51341.2" *)
  LUT4 \builder_count_mod_RNO_cZ[4]_TMR_0  (
    .A(N_699_TMR_0),
    .B(builder_wait_TMR_0),
    .C(sys_rst_TMR_0),
    .D(GND_0),
    .Z(builder_count_mod_RNO_TMR_0[4])
  );
  defparam \builder_count_mod_RNO_cZ[4]_TMR_0 .INIT = "0x0808";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51335.8-51341.2" *)
  LUT4 \builder_count_mod_RNO_cZ[4]_TMR_1  (
    .A(N_699_TMR_1),
    .B(builder_wait_TMR_1),
    .C(sys_rst_TMR_1),
    .D(GND_0),
    .Z(builder_count_mod_RNO_TMR_1[4])
  );
  defparam \builder_count_mod_RNO_cZ[4]_TMR_1 .INIT = "0x0808";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51335.8-51341.2" *)
  LUT4 \builder_count_mod_RNO_cZ[4]_TMR_2  (
    .A(N_699_TMR_2),
    .B(builder_wait_TMR_2),
    .C(sys_rst_TMR_2),
    .D(GND_0),
    .Z(builder_count_mod_RNO_TMR_2[4])
  );
  defparam \builder_count_mod_RNO_cZ[4]_TMR_2 .INIT = "0x0808";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51527.11-51538.2" *)
  WIDEFN9 \builder_csr_bankarray_dat_r_7_1_.m10_TMR_0  (
    .A0(m3_TMR_0),
    .A1(mem_adr0_TMR_0[0]),
    .B0(mem_adr0_TMR_0[0]),
    .B1(mem_adr0_TMR_0[1]),
    .C0(mem_adr0_TMR_0[2]),
    .C1(mem_adr0_TMR_0[2]),
    .D0(mem_adr0_TMR_0[3]),
    .D1(mem_adr0_TMR_0[3]),
    .SEL(mem_adr0_TMR_0[4]),
    .Z(m10_TMR_0)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m10_TMR_0 .INIT0 = "0xc355";
  defparam \builder_csr_bankarray_dat_r_7_1_.m10_TMR_0 .INIT1 = "0xd46b";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51527.11-51538.2" *)
  WIDEFN9 \builder_csr_bankarray_dat_r_7_1_.m10_TMR_1  (
    .A0(m3_TMR_1),
    .A1(mem_adr0_TMR_1[0]),
    .B0(mem_adr0_TMR_1[0]),
    .B1(mem_adr0_TMR_1[1]),
    .C0(mem_adr0_TMR_1[2]),
    .C1(mem_adr0_TMR_1[2]),
    .D0(mem_adr0_TMR_1[3]),
    .D1(mem_adr0_TMR_1[3]),
    .SEL(mem_adr0_TMR_1[4]),
    .Z(m10_TMR_1)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m10_TMR_1 .INIT0 = "0xc355";
  defparam \builder_csr_bankarray_dat_r_7_1_.m10_TMR_1 .INIT1 = "0xd46b";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51527.11-51538.2" *)
  WIDEFN9 \builder_csr_bankarray_dat_r_7_1_.m10_TMR_2  (
    .A0(m3_TMR_2),
    .A1(mem_adr0_TMR_2[0]),
    .B0(mem_adr0_TMR_2[0]),
    .B1(mem_adr0_TMR_2[1]),
    .C0(mem_adr0_TMR_2[2]),
    .C1(mem_adr0_TMR_2[2]),
    .D0(mem_adr0_TMR_2[3]),
    .D1(mem_adr0_TMR_2[3]),
    .SEL(mem_adr0_TMR_2[4]),
    .Z(m10_TMR_2)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m10_TMR_2 .INIT0 = "0xc355";
  defparam \builder_csr_bankarray_dat_r_7_1_.m10_TMR_2 .INIT1 = "0xd46b";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55996.8-56002.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m11_TMR_0  (
    .A(mem_adr0_TMR_0[0]),
    .B(mem_adr0_TMR_0[1]),
    .C(mem_adr0_TMR_0[2]),
    .D(GND_0),
    .Z(m11_TMR_0)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m11_TMR_0 .INIT = "0x3939";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55996.8-56002.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m11_TMR_1  (
    .A(mem_adr0_TMR_1[0]),
    .B(mem_adr0_TMR_1[1]),
    .C(mem_adr0_TMR_1[2]),
    .D(GND_0),
    .Z(m11_TMR_1)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m11_TMR_1 .INIT = "0x3939";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55996.8-56002.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m11_TMR_2  (
    .A(mem_adr0_TMR_2[0]),
    .B(mem_adr0_TMR_2[1]),
    .C(mem_adr0_TMR_2[2]),
    .D(GND_0),
    .Z(m11_TMR_2)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m11_TMR_2 .INIT = "0x3939";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56228.8-56234.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m12_TMR_0  (
    .A(mem_adr0_TMR_0[0]),
    .B(mem_adr0_TMR_0[2]),
    .C(GND_0),
    .D(GND_0),
    .Z(\builder_csr_bankarray_dat_r_7_1_.N_13_i_TMR_0 )
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m12_TMR_0 .INIT = "0x8888";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56228.8-56234.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m12_TMR_1  (
    .A(mem_adr0_TMR_1[0]),
    .B(mem_adr0_TMR_1[2]),
    .C(GND_0),
    .D(GND_0),
    .Z(\builder_csr_bankarray_dat_r_7_1_.N_13_i_TMR_1 )
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m12_TMR_1 .INIT = "0x8888";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56228.8-56234.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m12_TMR_2  (
    .A(mem_adr0_TMR_2[0]),
    .B(mem_adr0_TMR_2[2]),
    .C(GND_0),
    .D(GND_0),
    .Z(\builder_csr_bankarray_dat_r_7_1_.N_13_i_TMR_2 )
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m12_TMR_2 .INIT = "0x8888";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51512.11-51523.2" *)
  WIDEFN9 \builder_csr_bankarray_dat_r_7_1_.m18_TMR_0  (
    .A0(mem_adr0_TMR_0[3]),
    .A1(mem_adr0_TMR_0[0]),
    .B0(m11_TMR_0),
    .B1(mem_adr0_TMR_0[1]),
    .C0(mem_adr0_TMR_0[2]),
    .C1(mem_adr0_TMR_0[2]),
    .D0(mem_adr0_TMR_0[0]),
    .D1(mem_adr0_TMR_0[3]),
    .SEL(mem_adr0_TMR_0[4]),
    .Z(m18_TMR_0)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m18_TMR_0 .INIT0 = "0x3111";
  defparam \builder_csr_bankarray_dat_r_7_1_.m18_TMR_0 .INIT1 = "0x06d6";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51512.11-51523.2" *)
  WIDEFN9 \builder_csr_bankarray_dat_r_7_1_.m18_TMR_1  (
    .A0(mem_adr0_TMR_1[3]),
    .A1(mem_adr0_TMR_1[0]),
    .B0(m11_TMR_1),
    .B1(mem_adr0_TMR_1[1]),
    .C0(mem_adr0_TMR_1[2]),
    .C1(mem_adr0_TMR_1[2]),
    .D0(mem_adr0_TMR_1[0]),
    .D1(mem_adr0_TMR_1[3]),
    .SEL(mem_adr0_TMR_1[4]),
    .Z(m18_TMR_1)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m18_TMR_1 .INIT0 = "0x3111";
  defparam \builder_csr_bankarray_dat_r_7_1_.m18_TMR_1 .INIT1 = "0x06d6";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51512.11-51523.2" *)
  WIDEFN9 \builder_csr_bankarray_dat_r_7_1_.m18_TMR_2  (
    .A0(mem_adr0_TMR_2[3]),
    .A1(mem_adr0_TMR_2[0]),
    .B0(m11_TMR_2),
    .B1(mem_adr0_TMR_2[1]),
    .C0(mem_adr0_TMR_2[2]),
    .C1(mem_adr0_TMR_2[2]),
    .D0(mem_adr0_TMR_2[0]),
    .D1(mem_adr0_TMR_2[3]),
    .SEL(mem_adr0_TMR_2[4]),
    .Z(m18_TMR_2)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m18_TMR_2 .INIT0 = "0x3111";
  defparam \builder_csr_bankarray_dat_r_7_1_.m18_TMR_2 .INIT1 = "0x06d6";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56273.8-56279.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m19_TMR_0  (
    .A(m10_TMR_0),
    .B(m18_TMR_0),
    .C(mem_adr0_TMR_0[5]),
    .D(GND_0),
    .Z(builder_csr_bankarray_dat_r_TMR_0[1])
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m19_TMR_0 .INIT = "0xCACA";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56273.8-56279.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m19_TMR_1  (
    .A(m10_TMR_1),
    .B(m18_TMR_1),
    .C(mem_adr0_TMR_1[5]),
    .D(GND_0),
    .Z(builder_csr_bankarray_dat_r_TMR_1[1])
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m19_TMR_1 .INIT = "0xCACA";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56273.8-56279.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m19_TMR_2  (
    .A(m10_TMR_2),
    .B(m18_TMR_2),
    .C(mem_adr0_TMR_2[5]),
    .D(GND_0),
    .Z(builder_csr_bankarray_dat_r_TMR_2[1])
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m19_TMR_2 .INIT = "0xCACA";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55897.8-55903.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m30_TMR_0  (
    .A(mem_adr0_TMR_0[0]),
    .B(mem_adr0_TMR_0[1]),
    .C(mem_adr0_TMR_0[2]),
    .D(mem_adr0_TMR_0[3]),
    .Z(m30_TMR_0)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m30_TMR_0 .INIT = "0x696C";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55897.8-55903.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m30_TMR_1  (
    .A(mem_adr0_TMR_1[0]),
    .B(mem_adr0_TMR_1[1]),
    .C(mem_adr0_TMR_1[2]),
    .D(mem_adr0_TMR_1[3]),
    .Z(m30_TMR_1)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m30_TMR_1 .INIT = "0x696C";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55897.8-55903.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m30_TMR_2  (
    .A(mem_adr0_TMR_2[0]),
    .B(mem_adr0_TMR_2[1]),
    .C(mem_adr0_TMR_2[2]),
    .D(mem_adr0_TMR_2[3]),
    .Z(m30_TMR_2)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m30_TMR_2 .INIT = "0x696C";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55888.8-55894.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m33_TMR_0  (
    .A(mem_adr0_TMR_0[0]),
    .B(mem_adr0_TMR_0[1]),
    .C(mem_adr0_TMR_0[2]),
    .D(mem_adr0_TMR_0[3]),
    .Z(\builder_csr_bankarray_dat_r_7_1_.i2_mux_0_TMR_0 )
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m33_TMR_0 .INIT = "0x3D1A";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55888.8-55894.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m33_TMR_1  (
    .A(mem_adr0_TMR_1[0]),
    .B(mem_adr0_TMR_1[1]),
    .C(mem_adr0_TMR_1[2]),
    .D(mem_adr0_TMR_1[3]),
    .Z(\builder_csr_bankarray_dat_r_7_1_.i2_mux_0_TMR_1 )
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m33_TMR_1 .INIT = "0x3D1A";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55888.8-55894.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m33_TMR_2  (
    .A(mem_adr0_TMR_2[0]),
    .B(mem_adr0_TMR_2[1]),
    .C(mem_adr0_TMR_2[2]),
    .D(mem_adr0_TMR_2[3]),
    .Z(\builder_csr_bankarray_dat_r_7_1_.i2_mux_0_TMR_2 )
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m33_TMR_2 .INIT = "0x3D1A";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51557.11-51568.2" *)
  WIDEFN9 \builder_csr_bankarray_dat_r_7_1_.m35_TMR_0  (
    .A0(\builder_csr_bankarray_dat_r_7_1_.m35_am_1_TMR_0 ),
    .A1(m30_TMR_0),
    .B0(mem_adr0_TMR_0[1]),
    .B1(\builder_csr_bankarray_dat_r_7_1_.i2_mux_0_TMR_0 ),
    .C0(mem_adr0_TMR_0[3]),
    .C1(mem_adr0_TMR_0[4]),
    .D0(mem_adr0_TMR_0[4]),
    .D1(GND_0),
    .SEL(mem_adr0_TMR_0[5]),
    .Z(builder_csr_bankarray_dat_r_TMR_0[2])
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m35_TMR_0 .INIT0 = "0x87d4";
  defparam \builder_csr_bankarray_dat_r_7_1_.m35_TMR_0 .INIT1 = "0xcaca";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51557.11-51568.2" *)
  WIDEFN9 \builder_csr_bankarray_dat_r_7_1_.m35_TMR_1  (
    .A0(\builder_csr_bankarray_dat_r_7_1_.m35_am_1_TMR_1 ),
    .A1(m30_TMR_1),
    .B0(mem_adr0_TMR_1[1]),
    .B1(\builder_csr_bankarray_dat_r_7_1_.i2_mux_0_TMR_1 ),
    .C0(mem_adr0_TMR_1[3]),
    .C1(mem_adr0_TMR_1[4]),
    .D0(mem_adr0_TMR_1[4]),
    .D1(GND_0),
    .SEL(mem_adr0_TMR_1[5]),
    .Z(builder_csr_bankarray_dat_r_TMR_1[2])
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m35_TMR_1 .INIT0 = "0x87d4";
  defparam \builder_csr_bankarray_dat_r_7_1_.m35_TMR_1 .INIT1 = "0xcaca";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51557.11-51568.2" *)
  WIDEFN9 \builder_csr_bankarray_dat_r_7_1_.m35_TMR_2  (
    .A0(\builder_csr_bankarray_dat_r_7_1_.m35_am_1_TMR_2 ),
    .A1(m30_TMR_2),
    .B0(mem_adr0_TMR_2[1]),
    .B1(\builder_csr_bankarray_dat_r_7_1_.i2_mux_0_TMR_2 ),
    .C0(mem_adr0_TMR_2[3]),
    .C1(mem_adr0_TMR_2[4]),
    .D0(mem_adr0_TMR_2[4]),
    .D1(GND_0),
    .SEL(mem_adr0_TMR_2[5]),
    .Z(builder_csr_bankarray_dat_r_TMR_2[2])
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m35_TMR_2 .INIT0 = "0x87d4";
  defparam \builder_csr_bankarray_dat_r_7_1_.m35_TMR_2 .INIT1 = "0xcaca";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56327.8-56333.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m35_am_1_cZ_TMR_0  (
    .A(mem_adr0_TMR_0[0]),
    .B(mem_adr0_TMR_0[2]),
    .C(mem_adr0_TMR_0[3]),
    .D(mem_adr0_TMR_0[4]),
    .Z(\builder_csr_bankarray_dat_r_7_1_.m35_am_1_TMR_0 )
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m35_am_1_cZ_TMR_0 .INIT = "0x2763";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56327.8-56333.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m35_am_1_cZ_TMR_1  (
    .A(mem_adr0_TMR_1[0]),
    .B(mem_adr0_TMR_1[2]),
    .C(mem_adr0_TMR_1[3]),
    .D(mem_adr0_TMR_1[4]),
    .Z(\builder_csr_bankarray_dat_r_7_1_.m35_am_1_TMR_1 )
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m35_am_1_cZ_TMR_1 .INIT = "0x2763";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56327.8-56333.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m35_am_1_cZ_TMR_2  (
    .A(mem_adr0_TMR_2[0]),
    .B(mem_adr0_TMR_2[2]),
    .C(mem_adr0_TMR_2[3]),
    .D(mem_adr0_TMR_2[4]),
    .Z(\builder_csr_bankarray_dat_r_7_1_.m35_am_1_TMR_2 )
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m35_am_1_cZ_TMR_2 .INIT = "0x2763";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55951.8-55957.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m3_TMR_0  (
    .A(mem_adr0_TMR_0[0]),
    .B(mem_adr0_TMR_0[1]),
    .C(mem_adr0_TMR_0[2]),
    .D(GND_0),
    .Z(m3_TMR_0)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m3_TMR_0 .INIT = "0x3535";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55951.8-55957.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m3_TMR_1  (
    .A(mem_adr0_TMR_1[0]),
    .B(mem_adr0_TMR_1[1]),
    .C(mem_adr0_TMR_1[2]),
    .D(GND_0),
    .Z(m3_TMR_1)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m3_TMR_1 .INIT = "0x3535";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55951.8-55957.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m3_TMR_2  (
    .A(mem_adr0_TMR_2[0]),
    .B(mem_adr0_TMR_2[1]),
    .C(mem_adr0_TMR_2[2]),
    .D(GND_0),
    .Z(m3_TMR_2)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m3_TMR_2 .INIT = "0x3535";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51497.11-51508.2" *)
  WIDEFN9 \builder_csr_bankarray_dat_r_7_1_.m40_TMR_0  (
    .A0(mem_adr0_TMR_0[0]),
    .A1(m8_TMR_0),
    .B0(mem_adr0_TMR_0[1]),
    .B1(\builder_csr_bankarray_dat_r_7_1_.N_13_i_TMR_0 ),
    .C0(mem_adr0_TMR_0[2]),
    .C1(mem_adr0_TMR_0[1]),
    .D0(mem_adr0_TMR_0[3]),
    .D1(mem_adr0_TMR_0[3]),
    .SEL(mem_adr0_TMR_0[4]),
    .Z(m40_TMR_0)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m40_TMR_0 .INIT0 = "0x8c8d";
  defparam \builder_csr_bankarray_dat_r_7_1_.m40_TMR_0 .INIT1 = "0x3c55";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51497.11-51508.2" *)
  WIDEFN9 \builder_csr_bankarray_dat_r_7_1_.m40_TMR_1  (
    .A0(mem_adr0_TMR_1[0]),
    .A1(m8_TMR_1),
    .B0(mem_adr0_TMR_1[1]),
    .B1(\builder_csr_bankarray_dat_r_7_1_.N_13_i_TMR_1 ),
    .C0(mem_adr0_TMR_1[2]),
    .C1(mem_adr0_TMR_1[1]),
    .D0(mem_adr0_TMR_1[3]),
    .D1(mem_adr0_TMR_1[3]),
    .SEL(mem_adr0_TMR_1[4]),
    .Z(m40_TMR_1)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m40_TMR_1 .INIT0 = "0x8c8d";
  defparam \builder_csr_bankarray_dat_r_7_1_.m40_TMR_1 .INIT1 = "0x3c55";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51497.11-51508.2" *)
  WIDEFN9 \builder_csr_bankarray_dat_r_7_1_.m40_TMR_2  (
    .A0(mem_adr0_TMR_2[0]),
    .A1(m8_TMR_2),
    .B0(mem_adr0_TMR_2[1]),
    .B1(\builder_csr_bankarray_dat_r_7_1_.N_13_i_TMR_2 ),
    .C0(mem_adr0_TMR_2[2]),
    .C1(mem_adr0_TMR_2[1]),
    .D0(mem_adr0_TMR_2[3]),
    .D1(mem_adr0_TMR_2[3]),
    .SEL(mem_adr0_TMR_2[4]),
    .Z(m40_TMR_2)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m40_TMR_2 .INIT0 = "0x8c8d";
  defparam \builder_csr_bankarray_dat_r_7_1_.m40_TMR_2 .INIT1 = "0x3c55";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55987.8-55993.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m41_TMR_0  (
    .A(mem_adr0_TMR_0[0]),
    .B(mem_adr0_TMR_0[2]),
    .C(mem_adr0_TMR_0[3]),
    .D(GND_0),
    .Z(\builder_csr_bankarray_dat_r_7_1_.i3_mux_3_TMR_0 )
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m41_TMR_0 .INIT = "0xDEDE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55987.8-55993.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m41_TMR_1  (
    .A(mem_adr0_TMR_1[0]),
    .B(mem_adr0_TMR_1[2]),
    .C(mem_adr0_TMR_1[3]),
    .D(GND_0),
    .Z(\builder_csr_bankarray_dat_r_7_1_.i3_mux_3_TMR_1 )
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m41_TMR_1 .INIT = "0xDEDE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55987.8-55993.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m41_TMR_2  (
    .A(mem_adr0_TMR_2[0]),
    .B(mem_adr0_TMR_2[2]),
    .C(mem_adr0_TMR_2[3]),
    .D(GND_0),
    .Z(\builder_csr_bankarray_dat_r_7_1_.i3_mux_3_TMR_2 )
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m41_TMR_2 .INIT = "0xDEDE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51482.11-51493.2" *)
  WIDEFN9 \builder_csr_bankarray_dat_r_7_1_.m45_TMR_0  (
    .A0(\builder_csr_bankarray_dat_r_7_1_.N_13_i_TMR_0 ),
    .A1(mem_adr0_TMR_0[0]),
    .B0(\builder_csr_bankarray_dat_r_7_1_.i3_mux_3_TMR_0 ),
    .B1(mem_adr0_TMR_0[1]),
    .C0(mem_adr0_TMR_0[1]),
    .C1(mem_adr0_TMR_0[2]),
    .D0(mem_adr0_TMR_0[3]),
    .D1(mem_adr0_TMR_0[3]),
    .SEL(mem_adr0_TMR_0[4]),
    .Z(m45_TMR_0)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m45_TMR_0 .INIT0 = "0xa353";
  defparam \builder_csr_bankarray_dat_r_7_1_.m45_TMR_0 .INIT1 = "0x0696";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51482.11-51493.2" *)
  WIDEFN9 \builder_csr_bankarray_dat_r_7_1_.m45_TMR_1  (
    .A0(\builder_csr_bankarray_dat_r_7_1_.N_13_i_TMR_1 ),
    .A1(mem_adr0_TMR_1[0]),
    .B0(\builder_csr_bankarray_dat_r_7_1_.i3_mux_3_TMR_1 ),
    .B1(mem_adr0_TMR_1[1]),
    .C0(mem_adr0_TMR_1[1]),
    .C1(mem_adr0_TMR_1[2]),
    .D0(mem_adr0_TMR_1[3]),
    .D1(mem_adr0_TMR_1[3]),
    .SEL(mem_adr0_TMR_1[4]),
    .Z(m45_TMR_1)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m45_TMR_1 .INIT0 = "0xa353";
  defparam \builder_csr_bankarray_dat_r_7_1_.m45_TMR_1 .INIT1 = "0x0696";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51482.11-51493.2" *)
  WIDEFN9 \builder_csr_bankarray_dat_r_7_1_.m45_TMR_2  (
    .A0(\builder_csr_bankarray_dat_r_7_1_.N_13_i_TMR_2 ),
    .A1(mem_adr0_TMR_2[0]),
    .B0(\builder_csr_bankarray_dat_r_7_1_.i3_mux_3_TMR_2 ),
    .B1(mem_adr0_TMR_2[1]),
    .C0(mem_adr0_TMR_2[1]),
    .C1(mem_adr0_TMR_2[2]),
    .D0(mem_adr0_TMR_2[3]),
    .D1(mem_adr0_TMR_2[3]),
    .SEL(mem_adr0_TMR_2[4]),
    .Z(m45_TMR_2)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m45_TMR_2 .INIT0 = "0xa353";
  defparam \builder_csr_bankarray_dat_r_7_1_.m45_TMR_2 .INIT1 = "0x0696";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56282.8-56288.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m46_TMR_0  (
    .A(m40_TMR_0),
    .B(m45_TMR_0),
    .C(mem_adr0_TMR_0[5]),
    .D(GND_0),
    .Z(builder_csr_bankarray_dat_r_TMR_0[3])
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m46_TMR_0 .INIT = "0xCACA";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56282.8-56288.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m46_TMR_1  (
    .A(m40_TMR_1),
    .B(m45_TMR_1),
    .C(mem_adr0_TMR_1[5]),
    .D(GND_0),
    .Z(builder_csr_bankarray_dat_r_TMR_1[3])
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m46_TMR_1 .INIT = "0xCACA";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56282.8-56288.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m46_TMR_2  (
    .A(m40_TMR_2),
    .B(m45_TMR_2),
    .C(mem_adr0_TMR_2[5]),
    .D(GND_0),
    .Z(builder_csr_bankarray_dat_r_TMR_2[3])
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m46_TMR_2 .INIT = "0xCACA";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51422.11-51433.2" *)
  WIDEFN9 \builder_csr_bankarray_dat_r_7_1_.m51_TMR_0  (
    .A0(m6_TMR_0),
    .A1(mem_adr0_TMR_0[0]),
    .B0(\builder_csr_bankarray_dat_r_7_1_.N_13_i_TMR_0 ),
    .B1(mem_adr0_TMR_0[1]),
    .C0(mem_adr0_TMR_0[1]),
    .C1(mem_adr0_TMR_0[2]),
    .D0(mem_adr0_TMR_0[3]),
    .D1(mem_adr0_TMR_0[3]),
    .SEL(mem_adr0_TMR_0[4]),
    .Z(m51_TMR_0)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m51_TMR_0 .INIT0 = "0x50c3";
  defparam \builder_csr_bankarray_dat_r_7_1_.m51_TMR_0 .INIT1 = "0x21fc";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51422.11-51433.2" *)
  WIDEFN9 \builder_csr_bankarray_dat_r_7_1_.m51_TMR_1  (
    .A0(m6_TMR_1),
    .A1(mem_adr0_TMR_1[0]),
    .B0(\builder_csr_bankarray_dat_r_7_1_.N_13_i_TMR_1 ),
    .B1(mem_adr0_TMR_1[1]),
    .C0(mem_adr0_TMR_1[1]),
    .C1(mem_adr0_TMR_1[2]),
    .D0(mem_adr0_TMR_1[3]),
    .D1(mem_adr0_TMR_1[3]),
    .SEL(mem_adr0_TMR_1[4]),
    .Z(m51_TMR_1)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m51_TMR_1 .INIT0 = "0x50c3";
  defparam \builder_csr_bankarray_dat_r_7_1_.m51_TMR_1 .INIT1 = "0x21fc";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51422.11-51433.2" *)
  WIDEFN9 \builder_csr_bankarray_dat_r_7_1_.m51_TMR_2  (
    .A0(m6_TMR_2),
    .A1(mem_adr0_TMR_2[0]),
    .B0(\builder_csr_bankarray_dat_r_7_1_.N_13_i_TMR_2 ),
    .B1(mem_adr0_TMR_2[1]),
    .C0(mem_adr0_TMR_2[1]),
    .C1(mem_adr0_TMR_2[2]),
    .D0(mem_adr0_TMR_2[3]),
    .D1(mem_adr0_TMR_2[3]),
    .SEL(mem_adr0_TMR_2[4]),
    .Z(m51_TMR_2)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m51_TMR_2 .INIT0 = "0x50c3";
  defparam \builder_csr_bankarray_dat_r_7_1_.m51_TMR_2 .INIT1 = "0x21fc";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55969.8-55975.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m52_TMR_0  (
    .A(mem_adr0_TMR_0[0]),
    .B(mem_adr0_TMR_0[1]),
    .C(mem_adr0_TMR_0[2]),
    .D(GND_0),
    .Z(m52_TMR_0)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m52_TMR_0 .INIT = "0x4E4E";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55969.8-55975.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m52_TMR_1  (
    .A(mem_adr0_TMR_1[0]),
    .B(mem_adr0_TMR_1[1]),
    .C(mem_adr0_TMR_1[2]),
    .D(GND_0),
    .Z(m52_TMR_1)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m52_TMR_1 .INIT = "0x4E4E";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55969.8-55975.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m52_TMR_2  (
    .A(mem_adr0_TMR_2[0]),
    .B(mem_adr0_TMR_2[1]),
    .C(mem_adr0_TMR_2[2]),
    .D(GND_0),
    .Z(m52_TMR_2)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m52_TMR_2 .INIT = "0x4E4E";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51467.11-51478.2" *)
  WIDEFN9 \builder_csr_bankarray_dat_r_7_1_.m57_TMR_0  (
    .A0(m52_TMR_0),
    .A1(mem_adr0_TMR_0[0]),
    .B0(mem_adr0_TMR_0[1]),
    .B1(mem_adr0_TMR_0[1]),
    .C0(mem_adr0_TMR_0[3]),
    .C1(mem_adr0_TMR_0[2]),
    .D0(GND_0),
    .D1(mem_adr0_TMR_0[3]),
    .SEL(mem_adr0_TMR_0[4]),
    .Z(m57_TMR_0)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m57_TMR_0 .INIT0 = "0x4a4a";
  defparam \builder_csr_bankarray_dat_r_7_1_.m57_TMR_0 .INIT1 = "0x0904";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51467.11-51478.2" *)
  WIDEFN9 \builder_csr_bankarray_dat_r_7_1_.m57_TMR_1  (
    .A0(m52_TMR_1),
    .A1(mem_adr0_TMR_1[0]),
    .B0(mem_adr0_TMR_1[1]),
    .B1(mem_adr0_TMR_1[1]),
    .C0(mem_adr0_TMR_1[3]),
    .C1(mem_adr0_TMR_1[2]),
    .D0(GND_0),
    .D1(mem_adr0_TMR_1[3]),
    .SEL(mem_adr0_TMR_1[4]),
    .Z(m57_TMR_1)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m57_TMR_1 .INIT0 = "0x4a4a";
  defparam \builder_csr_bankarray_dat_r_7_1_.m57_TMR_1 .INIT1 = "0x0904";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51467.11-51478.2" *)
  WIDEFN9 \builder_csr_bankarray_dat_r_7_1_.m57_TMR_2  (
    .A0(m52_TMR_2),
    .A1(mem_adr0_TMR_2[0]),
    .B0(mem_adr0_TMR_2[1]),
    .B1(mem_adr0_TMR_2[1]),
    .C0(mem_adr0_TMR_2[3]),
    .C1(mem_adr0_TMR_2[2]),
    .D0(GND_0),
    .D1(mem_adr0_TMR_2[3]),
    .SEL(mem_adr0_TMR_2[4]),
    .Z(m57_TMR_2)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m57_TMR_2 .INIT0 = "0x4a4a";
  defparam \builder_csr_bankarray_dat_r_7_1_.m57_TMR_2 .INIT1 = "0x0904";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56291.8-56297.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m58_TMR_0  (
    .A(m51_TMR_0),
    .B(m57_TMR_0),
    .C(mem_adr0_TMR_0[5]),
    .D(GND_0),
    .Z(builder_csr_bankarray_dat_r_TMR_0[4])
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m58_TMR_0 .INIT = "0xCACA";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56291.8-56297.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m58_TMR_1  (
    .A(m51_TMR_1),
    .B(m57_TMR_1),
    .C(mem_adr0_TMR_1[5]),
    .D(GND_0),
    .Z(builder_csr_bankarray_dat_r_TMR_1[4])
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m58_TMR_1 .INIT = "0xCACA";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56291.8-56297.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m58_TMR_2  (
    .A(m51_TMR_2),
    .B(m57_TMR_2),
    .C(mem_adr0_TMR_2[5]),
    .D(GND_0),
    .Z(builder_csr_bankarray_dat_r_TMR_2[4])
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m58_TMR_2 .INIT = "0xCACA";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51452.11-51463.2" *)
  WIDEFN9 \builder_csr_bankarray_dat_r_7_1_.m64_TMR_0  (
    .A0(m6_TMR_0),
    .A1(mem_adr0_TMR_0[0]),
    .B0(mem_adr0_TMR_0[0]),
    .B1(mem_adr0_TMR_0[1]),
    .C0(mem_adr0_TMR_0[1]),
    .C1(mem_adr0_TMR_0[2]),
    .D0(mem_adr0_TMR_0[3]),
    .D1(mem_adr0_TMR_0[3]),
    .SEL(mem_adr0_TMR_0[4]),
    .Z(m64_TMR_0)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m64_TMR_0 .INIT0 = "0x5fc5";
  defparam \builder_csr_bankarray_dat_r_7_1_.m64_TMR_0 .INIT1 = "0xb6fc";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51452.11-51463.2" *)
  WIDEFN9 \builder_csr_bankarray_dat_r_7_1_.m64_TMR_1  (
    .A0(m6_TMR_1),
    .A1(mem_adr0_TMR_1[0]),
    .B0(mem_adr0_TMR_1[0]),
    .B1(mem_adr0_TMR_1[1]),
    .C0(mem_adr0_TMR_1[1]),
    .C1(mem_adr0_TMR_1[2]),
    .D0(mem_adr0_TMR_1[3]),
    .D1(mem_adr0_TMR_1[3]),
    .SEL(mem_adr0_TMR_1[4]),
    .Z(m64_TMR_1)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m64_TMR_1 .INIT0 = "0x5fc5";
  defparam \builder_csr_bankarray_dat_r_7_1_.m64_TMR_1 .INIT1 = "0xb6fc";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51452.11-51463.2" *)
  WIDEFN9 \builder_csr_bankarray_dat_r_7_1_.m64_TMR_2  (
    .A0(m6_TMR_2),
    .A1(mem_adr0_TMR_2[0]),
    .B0(mem_adr0_TMR_2[0]),
    .B1(mem_adr0_TMR_2[1]),
    .C0(mem_adr0_TMR_2[1]),
    .C1(mem_adr0_TMR_2[2]),
    .D0(mem_adr0_TMR_2[3]),
    .D1(mem_adr0_TMR_2[3]),
    .SEL(mem_adr0_TMR_2[4]),
    .Z(m64_TMR_2)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m64_TMR_2 .INIT0 = "0x5fc5";
  defparam \builder_csr_bankarray_dat_r_7_1_.m64_TMR_2 .INIT1 = "0xb6fc";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55978.8-55984.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m68_TMR_0  (
    .A(mem_adr0_TMR_0[0]),
    .B(mem_adr0_TMR_0[1]),
    .C(mem_adr0_TMR_0[2]),
    .D(GND_0),
    .Z(m68_TMR_0)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m68_TMR_0 .INIT = "0x2424";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55978.8-55984.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m68_TMR_1  (
    .A(mem_adr0_TMR_1[0]),
    .B(mem_adr0_TMR_1[1]),
    .C(mem_adr0_TMR_1[2]),
    .D(GND_0),
    .Z(m68_TMR_1)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m68_TMR_1 .INIT = "0x2424";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55978.8-55984.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m68_TMR_2  (
    .A(mem_adr0_TMR_2[0]),
    .B(mem_adr0_TMR_2[1]),
    .C(mem_adr0_TMR_2[2]),
    .D(GND_0),
    .Z(m68_TMR_2)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m68_TMR_2 .INIT = "0x2424";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56219.8-56225.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m6_TMR_0  (
    .A(mem_adr0_TMR_0[0]),
    .B(mem_adr0_TMR_0[2]),
    .C(GND_0),
    .D(GND_0),
    .Z(m6_TMR_0)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m6_TMR_0 .INIT = "0x4444";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56219.8-56225.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m6_TMR_1  (
    .A(mem_adr0_TMR_1[0]),
    .B(mem_adr0_TMR_1[2]),
    .C(GND_0),
    .D(GND_0),
    .Z(m6_TMR_1)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m6_TMR_1 .INIT = "0x4444";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56219.8-56225.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m6_TMR_2  (
    .A(mem_adr0_TMR_2[0]),
    .B(mem_adr0_TMR_2[2]),
    .C(GND_0),
    .D(GND_0),
    .Z(m6_TMR_2)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m6_TMR_2 .INIT = "0x4444";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51437.11-51448.2" *)
  WIDEFN9 \builder_csr_bankarray_dat_r_7_1_.m70_TMR_0  (
    .A0(mem_adr0_TMR_0[0]),
    .A1(m6_TMR_0),
    .B0(mem_adr0_TMR_0[1]),
    .B1(m68_TMR_0),
    .C0(mem_adr0_TMR_0[2]),
    .C1(mem_adr0_TMR_0[1]),
    .D0(mem_adr0_TMR_0[3]),
    .D1(mem_adr0_TMR_0[3]),
    .SEL(mem_adr0_TMR_0[4]),
    .Z(m70_TMR_0)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m70_TMR_0 .INIT0 = "0x86fe";
  defparam \builder_csr_bankarray_dat_r_7_1_.m70_TMR_0 .INIT1 = "0xa0cc";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51437.11-51448.2" *)
  WIDEFN9 \builder_csr_bankarray_dat_r_7_1_.m70_TMR_1  (
    .A0(mem_adr0_TMR_1[0]),
    .A1(m6_TMR_1),
    .B0(mem_adr0_TMR_1[1]),
    .B1(m68_TMR_1),
    .C0(mem_adr0_TMR_1[2]),
    .C1(mem_adr0_TMR_1[1]),
    .D0(mem_adr0_TMR_1[3]),
    .D1(mem_adr0_TMR_1[3]),
    .SEL(mem_adr0_TMR_1[4]),
    .Z(m70_TMR_1)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m70_TMR_1 .INIT0 = "0x86fe";
  defparam \builder_csr_bankarray_dat_r_7_1_.m70_TMR_1 .INIT1 = "0xa0cc";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51437.11-51448.2" *)
  WIDEFN9 \builder_csr_bankarray_dat_r_7_1_.m70_TMR_2  (
    .A0(mem_adr0_TMR_2[0]),
    .A1(m6_TMR_2),
    .B0(mem_adr0_TMR_2[1]),
    .B1(m68_TMR_2),
    .C0(mem_adr0_TMR_2[2]),
    .C1(mem_adr0_TMR_2[1]),
    .D0(mem_adr0_TMR_2[3]),
    .D1(mem_adr0_TMR_2[3]),
    .SEL(mem_adr0_TMR_2[4]),
    .Z(m70_TMR_2)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m70_TMR_2 .INIT0 = "0x86fe";
  defparam \builder_csr_bankarray_dat_r_7_1_.m70_TMR_2 .INIT1 = "0xa0cc";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56300.8-56306.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m71_TMR_0  (
    .A(m64_TMR_0),
    .B(m70_TMR_0),
    .C(mem_adr0_TMR_0[5]),
    .D(GND_0),
    .Z(m71_TMR_0)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m71_TMR_0 .INIT = "0xCACA";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56300.8-56306.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m71_TMR_1  (
    .A(m64_TMR_1),
    .B(m70_TMR_1),
    .C(mem_adr0_TMR_1[5]),
    .D(GND_0),
    .Z(m71_TMR_1)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m71_TMR_1 .INIT = "0xCACA";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56300.8-56306.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m71_TMR_2  (
    .A(m64_TMR_2),
    .B(m70_TMR_2),
    .C(mem_adr0_TMR_2[5]),
    .D(GND_0),
    .Z(m71_TMR_2)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m71_TMR_2 .INIT = "0xCACA";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55879.8-55885.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m73_TMR_0  (
    .A(mem_adr0_TMR_0[0]),
    .B(mem_adr0_TMR_0[1]),
    .C(mem_adr0_TMR_0[2]),
    .D(mem_adr0_TMR_0[3]),
    .Z(m73_TMR_0)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m73_TMR_0 .INIT = "0x2151";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55879.8-55885.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m73_TMR_1  (
    .A(mem_adr0_TMR_1[0]),
    .B(mem_adr0_TMR_1[1]),
    .C(mem_adr0_TMR_1[2]),
    .D(mem_adr0_TMR_1[3]),
    .Z(m73_TMR_1)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m73_TMR_1 .INIT = "0x2151";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55879.8-55885.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m73_TMR_2  (
    .A(mem_adr0_TMR_2[0]),
    .B(mem_adr0_TMR_2[1]),
    .C(mem_adr0_TMR_2[2]),
    .D(mem_adr0_TMR_2[3]),
    .Z(m73_TMR_2)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m73_TMR_2 .INIT = "0x2151";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55906.8-55912.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m74_TMR_0  (
    .A(mem_adr0_TMR_0[0]),
    .B(mem_adr0_TMR_0[1]),
    .C(mem_adr0_TMR_0[2]),
    .D(mem_adr0_TMR_0[3]),
    .Z(m74_TMR_0)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m74_TMR_0 .INIT = "0x0580";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55906.8-55912.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m74_TMR_1  (
    .A(mem_adr0_TMR_1[0]),
    .B(mem_adr0_TMR_1[1]),
    .C(mem_adr0_TMR_1[2]),
    .D(mem_adr0_TMR_1[3]),
    .Z(m74_TMR_1)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m74_TMR_1 .INIT = "0x0580";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55906.8-55912.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m74_TMR_2  (
    .A(mem_adr0_TMR_2[0]),
    .B(mem_adr0_TMR_2[1]),
    .C(mem_adr0_TMR_2[2]),
    .D(mem_adr0_TMR_2[3]),
    .Z(m74_TMR_2)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m74_TMR_2 .INIT = "0x0580";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56344.8-56350.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m77_TMR_0  (
    .A(mem_adr0_TMR_0[4]),
    .B(mem_adr0_TMR_0[2]),
    .C(mem_adr0_TMR_0[1]),
    .D(mem_adr0_TMR_0[0]),
    .Z(\builder_csr_bankarray_dat_r_7_1_.i4_mux_TMR_0 )
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m77_TMR_0 .INIT = "0x7B7F";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56344.8-56350.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m77_TMR_1  (
    .A(mem_adr0_TMR_1[4]),
    .B(mem_adr0_TMR_1[2]),
    .C(mem_adr0_TMR_1[1]),
    .D(mem_adr0_TMR_1[0]),
    .Z(\builder_csr_bankarray_dat_r_7_1_.i4_mux_TMR_1 )
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m77_TMR_1 .INIT = "0x7B7F";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56344.8-56350.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m77_TMR_2  (
    .A(mem_adr0_TMR_2[4]),
    .B(mem_adr0_TMR_2[2]),
    .C(mem_adr0_TMR_2[1]),
    .D(mem_adr0_TMR_2[0]),
    .Z(\builder_csr_bankarray_dat_r_7_1_.i4_mux_TMR_2 )
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m77_TMR_2 .INIT = "0x7B7F";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51542.11-51553.2" *)
  WIDEFN9 \builder_csr_bankarray_dat_r_7_1_.m80_TMR_0  (
    .A0(m73_TMR_0),
    .A1(\builder_csr_bankarray_dat_r_7_1_.i4_mux_TMR_0 ),
    .B0(m74_TMR_0),
    .B1(mem_adr0_TMR_0[3]),
    .C0(mem_adr0_TMR_0[4]),
    .C1(mem_adr0_TMR_0[4]),
    .D0(GND_0),
    .D1(GND_0),
    .SEL(mem_adr0_TMR_0[5]),
    .Z(builder_csr_bankarray_dat_r_TMR_0[6])
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m80_TMR_0 .INIT0 = "0x3535";
  defparam \builder_csr_bankarray_dat_r_7_1_.m80_TMR_0 .INIT1 = "0xbebe";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51542.11-51553.2" *)
  WIDEFN9 \builder_csr_bankarray_dat_r_7_1_.m80_TMR_1  (
    .A0(m73_TMR_1),
    .A1(\builder_csr_bankarray_dat_r_7_1_.i4_mux_TMR_1 ),
    .B0(m74_TMR_1),
    .B1(mem_adr0_TMR_1[3]),
    .C0(mem_adr0_TMR_1[4]),
    .C1(mem_adr0_TMR_1[4]),
    .D0(GND_0),
    .D1(GND_0),
    .SEL(mem_adr0_TMR_1[5]),
    .Z(builder_csr_bankarray_dat_r_TMR_1[6])
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m80_TMR_1 .INIT0 = "0x3535";
  defparam \builder_csr_bankarray_dat_r_7_1_.m80_TMR_1 .INIT1 = "0xbebe";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51542.11-51553.2" *)
  WIDEFN9 \builder_csr_bankarray_dat_r_7_1_.m80_TMR_2  (
    .A0(m73_TMR_2),
    .A1(\builder_csr_bankarray_dat_r_7_1_.i4_mux_TMR_2 ),
    .B0(m74_TMR_2),
    .B1(mem_adr0_TMR_2[3]),
    .C0(mem_adr0_TMR_2[4]),
    .C1(mem_adr0_TMR_2[4]),
    .D0(GND_0),
    .D1(GND_0),
    .SEL(mem_adr0_TMR_2[5]),
    .Z(builder_csr_bankarray_dat_r_TMR_2[6])
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m80_TMR_2 .INIT0 = "0x3535";
  defparam \builder_csr_bankarray_dat_r_7_1_.m80_TMR_2 .INIT1 = "0xbebe";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51407.11-51418.2" *)
  WIDEFN9 \builder_csr_bankarray_dat_r_7_1_.m84_TMR_0  (
    .A0(mem_adr0_TMR_0[0]),
    .A1(mem_adr0_TMR_0[0]),
    .B0(mem_adr0_TMR_0[1]),
    .B1(mem_adr0_TMR_0[1]),
    .C0(mem_adr0_TMR_0[2]),
    .C1(mem_adr0_TMR_0[2]),
    .D0(mem_adr0_TMR_0[3]),
    .D1(mem_adr0_TMR_0[3]),
    .SEL(mem_adr0_TMR_0[4]),
    .Z(m84_TMR_0)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m84_TMR_0 .INIT0 = "0x1220";
  defparam \builder_csr_bankarray_dat_r_7_1_.m84_TMR_0 .INIT1 = "0x0240";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51407.11-51418.2" *)
  WIDEFN9 \builder_csr_bankarray_dat_r_7_1_.m84_TMR_1  (
    .A0(mem_adr0_TMR_1[0]),
    .A1(mem_adr0_TMR_1[0]),
    .B0(mem_adr0_TMR_1[1]),
    .B1(mem_adr0_TMR_1[1]),
    .C0(mem_adr0_TMR_1[2]),
    .C1(mem_adr0_TMR_1[2]),
    .D0(mem_adr0_TMR_1[3]),
    .D1(mem_adr0_TMR_1[3]),
    .SEL(mem_adr0_TMR_1[4]),
    .Z(m84_TMR_1)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m84_TMR_1 .INIT0 = "0x1220";
  defparam \builder_csr_bankarray_dat_r_7_1_.m84_TMR_1 .INIT1 = "0x0240";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51407.11-51418.2" *)
  WIDEFN9 \builder_csr_bankarray_dat_r_7_1_.m84_TMR_2  (
    .A0(mem_adr0_TMR_2[0]),
    .A1(mem_adr0_TMR_2[0]),
    .B0(mem_adr0_TMR_2[1]),
    .B1(mem_adr0_TMR_2[1]),
    .C0(mem_adr0_TMR_2[2]),
    .C1(mem_adr0_TMR_2[2]),
    .D0(mem_adr0_TMR_2[3]),
    .D1(mem_adr0_TMR_2[3]),
    .SEL(mem_adr0_TMR_2[4]),
    .Z(m84_TMR_2)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m84_TMR_2 .INIT0 = "0x1220";
  defparam \builder_csr_bankarray_dat_r_7_1_.m84_TMR_2 .INIT1 = "0x0240";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51353.8-51359.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m86_TMR_0  (
    .A(mem_adr0_TMR_0[3]),
    .B(mem_adr0_TMR_0[2]),
    .C(mem_adr0_TMR_0[1]),
    .D(mem_adr0_TMR_0[0]),
    .Z(m86_TMR_0)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m86_TMR_0 .INIT = "0x5753";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51353.8-51359.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m86_TMR_1  (
    .A(mem_adr0_TMR_1[3]),
    .B(mem_adr0_TMR_1[2]),
    .C(mem_adr0_TMR_1[1]),
    .D(mem_adr0_TMR_1[0]),
    .Z(m86_TMR_1)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m86_TMR_1 .INIT = "0x5753";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51353.8-51359.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m86_TMR_2  (
    .A(mem_adr0_TMR_2[3]),
    .B(mem_adr0_TMR_2[2]),
    .C(mem_adr0_TMR_2[1]),
    .D(mem_adr0_TMR_2[0]),
    .Z(m86_TMR_2)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m86_TMR_2 .INIT = "0x5753";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55800.8-55806.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m88_TMR_0  (
    .A(m84_TMR_0),
    .B(m86_TMR_0),
    .C(mem_adr0_TMR_0[4]),
    .D(mem_adr0_TMR_0[5]),
    .Z(builder_csr_bankarray_dat_r_TMR_0[7])
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m88_TMR_0 .INIT = "0x0C55";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55800.8-55806.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m88_TMR_1  (
    .A(m84_TMR_1),
    .B(m86_TMR_1),
    .C(mem_adr0_TMR_1[4]),
    .D(mem_adr0_TMR_1[5]),
    .Z(builder_csr_bankarray_dat_r_TMR_1[7])
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m88_TMR_1 .INIT = "0x0C55";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55800.8-55806.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m88_TMR_2  (
    .A(m84_TMR_2),
    .B(m86_TMR_2),
    .C(mem_adr0_TMR_2[4]),
    .D(mem_adr0_TMR_2[5]),
    .Z(builder_csr_bankarray_dat_r_TMR_2[7])
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m88_TMR_2 .INIT = "0x0C55";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55960.8-55966.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m8_TMR_0  (
    .A(mem_adr0_TMR_0[0]),
    .B(mem_adr0_TMR_0[1]),
    .C(mem_adr0_TMR_0[2]),
    .D(GND_0),
    .Z(m8_TMR_0)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m8_TMR_0 .INIT = "0x2B2B";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55960.8-55966.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m8_TMR_1  (
    .A(mem_adr0_TMR_1[0]),
    .B(mem_adr0_TMR_1[1]),
    .C(mem_adr0_TMR_1[2]),
    .D(GND_0),
    .Z(m8_TMR_1)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m8_TMR_1 .INIT = "0x2B2B";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55960.8-55966.2" *)
  LUT4 \builder_csr_bankarray_dat_r_7_1_.m8_TMR_2  (
    .A(mem_adr0_TMR_2[0]),
    .B(mem_adr0_TMR_2[1]),
    .C(mem_adr0_TMR_2[2]),
    .D(GND_0),
    .Z(m8_TMR_2)
  );
  defparam \builder_csr_bankarray_dat_r_7_1_.m8_TMR_2 .INIT = "0x2B2B";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55114.11-55120.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[0]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_0[0]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_0[0]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55114.11-55120.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[0]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_1[0]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_1[0]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55114.11-55120.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[0]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_2[0]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_2[0]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55177.11-55183.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[10]_TMR_0  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_0 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_0[10]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_0[10]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55177.11-55183.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[10]_TMR_1  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_1 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_1[10]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_1[10]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55177.11-55183.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[10]_TMR_2  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_2 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_2[10]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_2[10]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55184.11-55190.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[11]_TMR_0  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_0 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_0[11]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_0[11]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55184.11-55190.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[11]_TMR_1  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_1 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_1[11]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_1[11]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55184.11-55190.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[11]_TMR_2  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_2 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_2[11]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_2[11]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55191.11-55197.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[12]_TMR_0  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_0 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_0[12]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_0[12]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55191.11-55197.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[12]_TMR_1  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_1 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_1[12]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_1[12]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55191.11-55197.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[12]_TMR_2  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_2 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_2[12]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_2[12]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55198.11-55204.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[13]_TMR_0  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_0 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_0[13]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_0[13]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55198.11-55204.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[13]_TMR_1  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_1 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_1[13]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_1[13]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55198.11-55204.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[13]_TMR_2  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_2 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_2[13]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_2[13]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55205.11-55211.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[14]_TMR_0  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_0 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_0[14]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_0[14]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55205.11-55211.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[14]_TMR_1  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_1 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_1[14]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_1[14]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55205.11-55211.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[14]_TMR_2  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_2 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_2[14]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_2[14]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55212.11-55218.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[15]_TMR_0  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_0 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_0[15]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_0[15]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55212.11-55218.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[15]_TMR_1  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_1 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_1[15]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_1[15]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55212.11-55218.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[15]_TMR_2  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_2 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_2[15]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_2[15]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55219.11-55225.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[16]_TMR_0  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_0 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_0[16]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_0[16]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55219.11-55225.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[16]_TMR_1  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_1 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_1[16]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_1[16]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55219.11-55225.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[16]_TMR_2  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_2 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_2[16]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_2[16]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55226.11-55232.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[17]_TMR_0  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_0 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_0[17]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_0[17]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55226.11-55232.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[17]_TMR_1  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_1 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_1[17]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_1[17]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55226.11-55232.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[17]_TMR_2  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_2 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_2[17]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_2[17]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55233.11-55239.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[18]_TMR_0  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_0 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_0[18]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_0[18]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55233.11-55239.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[18]_TMR_1  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_1 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_1[18]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_1[18]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55233.11-55239.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[18]_TMR_2  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_2 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_2[18]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_2[18]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55240.11-55246.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[19]_TMR_0  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_0 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_0[19]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_0[19]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55240.11-55246.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[19]_TMR_1  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_1 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_1[19]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_1[19]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55240.11-55246.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[19]_TMR_2  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_2 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_2[19]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_2[19]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55247.11-55253.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[20]_TMR_0  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_0 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_0[20]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_0[20]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55247.11-55253.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[20]_TMR_1  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_1 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_1[20]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_1[20]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55247.11-55253.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[20]_TMR_2  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_2 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_2[20]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_2[20]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55254.11-55260.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[21]_TMR_0  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_0 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_0[21]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_0[21]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55254.11-55260.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[21]_TMR_1  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_1 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_1[21]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_1[21]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55254.11-55260.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[21]_TMR_2  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_2 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_2[21]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_2[21]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55261.11-55267.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[22]_TMR_0  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_0 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_0[22]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_0[22]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55261.11-55267.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[22]_TMR_1  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_1 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_1[22]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_1[22]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55261.11-55267.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[22]_TMR_2  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_2 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_2[22]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_2[22]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55268.11-55274.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[23]_TMR_0  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_0 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_0[23]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_0[23]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55268.11-55274.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[23]_TMR_1  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_1 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_1[23]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_1[23]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55268.11-55274.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[23]_TMR_2  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_2 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_2[23]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_2[23]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55275.11-55281.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[24]_TMR_0  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_0 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_0[24]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_0[24]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55275.11-55281.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[24]_TMR_1  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_1 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_1[24]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_1[24]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55275.11-55281.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[24]_TMR_2  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_2 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_2[24]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_2[24]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55282.11-55288.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[25]_TMR_0  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_0 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_0[25]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_0[25]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55282.11-55288.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[25]_TMR_1  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_1 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_1[25]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_1[25]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55282.11-55288.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[25]_TMR_2  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_2 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_2[25]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_2[25]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55289.11-55295.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[26]_TMR_0  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_0 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_0[26]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_0[26]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55289.11-55295.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[26]_TMR_1  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_1 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_1[26]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_1[26]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55289.11-55295.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[26]_TMR_2  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_2 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_2[26]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_2[26]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55296.11-55302.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[27]_TMR_0  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_0 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_0[27]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_0[27]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55296.11-55302.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[27]_TMR_1  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_1 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_1[27]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_1[27]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55296.11-55302.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[27]_TMR_2  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_2 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_2[27]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_2[27]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55303.11-55309.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[28]_TMR_0  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_0 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_0[28]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_0[28]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55303.11-55309.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[28]_TMR_1  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_1 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_1[28]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_1[28]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55303.11-55309.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[28]_TMR_2  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_2 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_2[28]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_2[28]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55310.11-55316.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[29]_TMR_0  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_0 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_0[29]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_0[29]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55310.11-55316.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[29]_TMR_1  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_1 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_1[29]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_1[29]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55310.11-55316.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[29]_TMR_2  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_2 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_2[29]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_2[29]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55121.11-55127.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[2]_TMR_0  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_0 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_0[2]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_0[2]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55121.11-55127.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[2]_TMR_1  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_1 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_1[2]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_1[2]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55121.11-55127.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[2]_TMR_2  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_2 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_2[2]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_2[2]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55317.11-55323.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[30]_TMR_0  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_0 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_0[30]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_0[30]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55317.11-55323.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[30]_TMR_1  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_1 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_1[30]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_1[30]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55317.11-55323.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[30]_TMR_2  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_2 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_2[30]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_2[30]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55324.11-55330.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[31]_TMR_0  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_0 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_0[31]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_0[31]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55324.11-55330.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[31]_TMR_1  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_1 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_1[31]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_1[31]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55324.11-55330.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[31]_TMR_2  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_2 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_2[31]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_2[31]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55128.11-55134.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[3]_TMR_0  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_0 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_0[3]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_0[3]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55128.11-55134.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[3]_TMR_1  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_1 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_1[3]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_1[3]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55128.11-55134.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[3]_TMR_2  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_2 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_2[3]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_2[3]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55135.11-55141.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[4]_TMR_0  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_0 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_0[4]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_0[4]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55135.11-55141.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[4]_TMR_1  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_1 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_1[4]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_1[4]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55135.11-55141.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[4]_TMR_2  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_2 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_2[4]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_2[4]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55142.11-55148.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[5]_TMR_0  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_0 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_0[5]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_0[5]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55142.11-55148.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[5]_TMR_1  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_1 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_1[5]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_1[5]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55142.11-55148.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[5]_TMR_2  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_2 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_2[5]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_2[5]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55149.11-55155.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[6]_TMR_0  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_0 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_0[6]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_0[6]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55149.11-55155.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[6]_TMR_1  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_1 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_1[6]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_1[6]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55149.11-55155.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[6]_TMR_2  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_2 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_2[6]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_2[6]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55156.11-55162.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[7]_TMR_0  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_0 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_0[7]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_0[7]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55156.11-55162.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[7]_TMR_1  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_1 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_1[7]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_1[7]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55156.11-55162.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[7]_TMR_2  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_2 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_2[7]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_2[7]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55163.11-55169.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[8]_TMR_0  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_0 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_0[8]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_0[8]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55163.11-55169.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[8]_TMR_1  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_1 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_1[8]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_1[8]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55163.11-55169.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[8]_TMR_2  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_2 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_2[8]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_2[8]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55170.11-55176.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[9]_TMR_0  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_0 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_0[9]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_0[9]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55170.11-55176.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[9]_TMR_1  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_1 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_1[9]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_1[9]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55170.11-55176.2" *)
  FD1P3IX \builder_csr_bankarray_interface0_bank_bus_dat_r_reg[9]_TMR_2  (
    .CD(\VexRiscv.IBusCachedPlugin_cache.builder_csr_bankarray_interface0_bank_bus_dat_r_6_sn_m4_0_iso_TMR_2 ),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface0_bank_bus_dat_r_6_TMR_2[9]),
    .Q(builder_csr_bankarray_interface0_bank_bus_dat_r_TMR_2[9]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55016.11-55022.2" *)
  FD1P3IX \builder_csr_bankarray_interface1_bank_bus_dat_r_reg[0]_TMR_0  (
    .CD(builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_0),
    .CK(sys_clk),
    .D(main_storage_TMR_0[0]),
    .Q(builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_0[0]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55016.11-55022.2" *)
  FD1P3IX \builder_csr_bankarray_interface1_bank_bus_dat_r_reg[0]_TMR_1  (
    .CD(builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_1),
    .CK(sys_clk),
    .D(main_storage_TMR_1[0]),
    .Q(builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_1[0]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55016.11-55022.2" *)
  FD1P3IX \builder_csr_bankarray_interface1_bank_bus_dat_r_reg[0]_TMR_2  (
    .CD(builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_2),
    .CK(sys_clk),
    .D(main_storage_TMR_2[0]),
    .Q(builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_2[0]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55086.11-55092.2" *)
  FD1P3IX \builder_csr_bankarray_interface1_bank_bus_dat_r_reg[10]_TMR_0  (
    .CD(builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_0),
    .CK(sys_clk),
    .D(main_storage_TMR_0[10]),
    .Q(builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_0[10]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55086.11-55092.2" *)
  FD1P3IX \builder_csr_bankarray_interface1_bank_bus_dat_r_reg[10]_TMR_1  (
    .CD(builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_1),
    .CK(sys_clk),
    .D(main_storage_TMR_1[10]),
    .Q(builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_1[10]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55086.11-55092.2" *)
  FD1P3IX \builder_csr_bankarray_interface1_bank_bus_dat_r_reg[10]_TMR_2  (
    .CD(builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_2),
    .CK(sys_clk),
    .D(main_storage_TMR_2[10]),
    .Q(builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_2[10]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55093.11-55099.2" *)
  FD1P3IX \builder_csr_bankarray_interface1_bank_bus_dat_r_reg[11]_TMR_0  (
    .CD(builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_0),
    .CK(sys_clk),
    .D(main_storage_TMR_0[11]),
    .Q(builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_0[11]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55093.11-55099.2" *)
  FD1P3IX \builder_csr_bankarray_interface1_bank_bus_dat_r_reg[11]_TMR_1  (
    .CD(builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_1),
    .CK(sys_clk),
    .D(main_storage_TMR_1[11]),
    .Q(builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_1[11]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55093.11-55099.2" *)
  FD1P3IX \builder_csr_bankarray_interface1_bank_bus_dat_r_reg[11]_TMR_2  (
    .CD(builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_2),
    .CK(sys_clk),
    .D(main_storage_TMR_2[11]),
    .Q(builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_2[11]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55100.11-55106.2" *)
  FD1P3IX \builder_csr_bankarray_interface1_bank_bus_dat_r_reg[12]_TMR_0  (
    .CD(builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_0),
    .CK(sys_clk),
    .D(main_storage_TMR_0[12]),
    .Q(builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_0[12]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55100.11-55106.2" *)
  FD1P3IX \builder_csr_bankarray_interface1_bank_bus_dat_r_reg[12]_TMR_1  (
    .CD(builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_1),
    .CK(sys_clk),
    .D(main_storage_TMR_1[12]),
    .Q(builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_1[12]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55100.11-55106.2" *)
  FD1P3IX \builder_csr_bankarray_interface1_bank_bus_dat_r_reg[12]_TMR_2  (
    .CD(builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_2),
    .CK(sys_clk),
    .D(main_storage_TMR_2[12]),
    .Q(builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_2[12]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55107.11-55113.2" *)
  FD1P3IX \builder_csr_bankarray_interface1_bank_bus_dat_r_reg[13]_TMR_0  (
    .CD(builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_0),
    .CK(sys_clk),
    .D(main_storage_TMR_0[13]),
    .Q(builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_0[13]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55107.11-55113.2" *)
  FD1P3IX \builder_csr_bankarray_interface1_bank_bus_dat_r_reg[13]_TMR_1  (
    .CD(builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_1),
    .CK(sys_clk),
    .D(main_storage_TMR_1[13]),
    .Q(builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_1[13]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55107.11-55113.2" *)
  FD1P3IX \builder_csr_bankarray_interface1_bank_bus_dat_r_reg[13]_TMR_2  (
    .CD(builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_2),
    .CK(sys_clk),
    .D(main_storage_TMR_2[13]),
    .Q(builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_2[13]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55023.11-55029.2" *)
  FD1P3IX \builder_csr_bankarray_interface1_bank_bus_dat_r_reg[1]_TMR_0  (
    .CD(builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_0),
    .CK(sys_clk),
    .D(main_storage_TMR_0[1]),
    .Q(builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_0[1]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55023.11-55029.2" *)
  FD1P3IX \builder_csr_bankarray_interface1_bank_bus_dat_r_reg[1]_TMR_1  (
    .CD(builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_1),
    .CK(sys_clk),
    .D(main_storage_TMR_1[1]),
    .Q(builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_1[1]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55023.11-55029.2" *)
  FD1P3IX \builder_csr_bankarray_interface1_bank_bus_dat_r_reg[1]_TMR_2  (
    .CD(builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_2),
    .CK(sys_clk),
    .D(main_storage_TMR_2[1]),
    .Q(builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_2[1]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55030.11-55036.2" *)
  FD1P3IX \builder_csr_bankarray_interface1_bank_bus_dat_r_reg[2]_TMR_0  (
    .CD(builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_0),
    .CK(sys_clk),
    .D(main_storage_TMR_0[2]),
    .Q(builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_0[2]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55030.11-55036.2" *)
  FD1P3IX \builder_csr_bankarray_interface1_bank_bus_dat_r_reg[2]_TMR_1  (
    .CD(builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_1),
    .CK(sys_clk),
    .D(main_storage_TMR_1[2]),
    .Q(builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_1[2]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55030.11-55036.2" *)
  FD1P3IX \builder_csr_bankarray_interface1_bank_bus_dat_r_reg[2]_TMR_2  (
    .CD(builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_2),
    .CK(sys_clk),
    .D(main_storage_TMR_2[2]),
    .Q(builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_2[2]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55037.11-55043.2" *)
  FD1P3IX \builder_csr_bankarray_interface1_bank_bus_dat_r_reg[3]_TMR_0  (
    .CD(builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_0),
    .CK(sys_clk),
    .D(main_storage_TMR_0[3]),
    .Q(builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_0[3]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55037.11-55043.2" *)
  FD1P3IX \builder_csr_bankarray_interface1_bank_bus_dat_r_reg[3]_TMR_1  (
    .CD(builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_1),
    .CK(sys_clk),
    .D(main_storage_TMR_1[3]),
    .Q(builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_1[3]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55037.11-55043.2" *)
  FD1P3IX \builder_csr_bankarray_interface1_bank_bus_dat_r_reg[3]_TMR_2  (
    .CD(builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_2),
    .CK(sys_clk),
    .D(main_storage_TMR_2[3]),
    .Q(builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_2[3]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55044.11-55050.2" *)
  FD1P3IX \builder_csr_bankarray_interface1_bank_bus_dat_r_reg[4]_TMR_0  (
    .CD(builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_0),
    .CK(sys_clk),
    .D(main_storage_TMR_0[4]),
    .Q(builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_0[4]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55044.11-55050.2" *)
  FD1P3IX \builder_csr_bankarray_interface1_bank_bus_dat_r_reg[4]_TMR_1  (
    .CD(builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_1),
    .CK(sys_clk),
    .D(main_storage_TMR_1[4]),
    .Q(builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_1[4]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55044.11-55050.2" *)
  FD1P3IX \builder_csr_bankarray_interface1_bank_bus_dat_r_reg[4]_TMR_2  (
    .CD(builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_2),
    .CK(sys_clk),
    .D(main_storage_TMR_2[4]),
    .Q(builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_2[4]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55051.11-55057.2" *)
  FD1P3IX \builder_csr_bankarray_interface1_bank_bus_dat_r_reg[5]_TMR_0  (
    .CD(builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_0),
    .CK(sys_clk),
    .D(main_storage_TMR_0[5]),
    .Q(builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_0[5]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55051.11-55057.2" *)
  FD1P3IX \builder_csr_bankarray_interface1_bank_bus_dat_r_reg[5]_TMR_1  (
    .CD(builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_1),
    .CK(sys_clk),
    .D(main_storage_TMR_1[5]),
    .Q(builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_1[5]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55051.11-55057.2" *)
  FD1P3IX \builder_csr_bankarray_interface1_bank_bus_dat_r_reg[5]_TMR_2  (
    .CD(builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_2),
    .CK(sys_clk),
    .D(main_storage_TMR_2[5]),
    .Q(builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_2[5]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55058.11-55064.2" *)
  FD1P3IX \builder_csr_bankarray_interface1_bank_bus_dat_r_reg[6]_TMR_0  (
    .CD(builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_0),
    .CK(sys_clk),
    .D(main_storage_TMR_0[6]),
    .Q(builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_0[6]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55058.11-55064.2" *)
  FD1P3IX \builder_csr_bankarray_interface1_bank_bus_dat_r_reg[6]_TMR_1  (
    .CD(builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_1),
    .CK(sys_clk),
    .D(main_storage_TMR_1[6]),
    .Q(builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_1[6]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55058.11-55064.2" *)
  FD1P3IX \builder_csr_bankarray_interface1_bank_bus_dat_r_reg[6]_TMR_2  (
    .CD(builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_2),
    .CK(sys_clk),
    .D(main_storage_TMR_2[6]),
    .Q(builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_2[6]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55065.11-55071.2" *)
  FD1P3IX \builder_csr_bankarray_interface1_bank_bus_dat_r_reg[7]_TMR_0  (
    .CD(builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_0),
    .CK(sys_clk),
    .D(main_storage_TMR_0[7]),
    .Q(builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_0[7]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55065.11-55071.2" *)
  FD1P3IX \builder_csr_bankarray_interface1_bank_bus_dat_r_reg[7]_TMR_1  (
    .CD(builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_1),
    .CK(sys_clk),
    .D(main_storage_TMR_1[7]),
    .Q(builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_1[7]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55065.11-55071.2" *)
  FD1P3IX \builder_csr_bankarray_interface1_bank_bus_dat_r_reg[7]_TMR_2  (
    .CD(builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_2),
    .CK(sys_clk),
    .D(main_storage_TMR_2[7]),
    .Q(builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_2[7]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55072.11-55078.2" *)
  FD1P3IX \builder_csr_bankarray_interface1_bank_bus_dat_r_reg[8]_TMR_0  (
    .CD(builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_0),
    .CK(sys_clk),
    .D(main_storage_TMR_0[8]),
    .Q(builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_0[8]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55072.11-55078.2" *)
  FD1P3IX \builder_csr_bankarray_interface1_bank_bus_dat_r_reg[8]_TMR_1  (
    .CD(builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_1),
    .CK(sys_clk),
    .D(main_storage_TMR_1[8]),
    .Q(builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_1[8]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55072.11-55078.2" *)
  FD1P3IX \builder_csr_bankarray_interface1_bank_bus_dat_r_reg[8]_TMR_2  (
    .CD(builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_2),
    .CK(sys_clk),
    .D(main_storage_TMR_2[8]),
    .Q(builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_2[8]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55079.11-55085.2" *)
  FD1P3IX \builder_csr_bankarray_interface1_bank_bus_dat_r_reg[9]_TMR_0  (
    .CD(builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_0),
    .CK(sys_clk),
    .D(main_storage_TMR_0[9]),
    .Q(builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_0[9]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55079.11-55085.2" *)
  FD1P3IX \builder_csr_bankarray_interface1_bank_bus_dat_r_reg[9]_TMR_1  (
    .CD(builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_1),
    .CK(sys_clk),
    .D(main_storage_TMR_1[9]),
    .Q(builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_1[9]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55079.11-55085.2" *)
  FD1P3IX \builder_csr_bankarray_interface1_bank_bus_dat_r_reg[9]_TMR_2  (
    .CD(builder_csr_bankarray_interface1_bank_bus_dat_r_0_sqmuxa_i_TMR_2),
    .CK(sys_clk),
    .D(main_storage_TMR_2[9]),
    .Q(builder_csr_bankarray_interface1_bank_bus_dat_r_TMR_2[9]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54792.11-54798.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[0]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_0[0]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_0[0]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54792.11-54798.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[0]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_1[0]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_1[0]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54792.11-54798.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[0]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_2[0]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_2[0]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54862.11-54868.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[10]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_0[10]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_0[10]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54862.11-54868.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[10]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_1[10]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_1[10]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54862.11-54868.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[10]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_2[10]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_2[10]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54869.11-54875.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[11]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_0[11]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_0[11]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54869.11-54875.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[11]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_1[11]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_1[11]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54869.11-54875.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[11]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_2[11]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_2[11]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54876.11-54882.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[12]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_0[12]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_0[12]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54876.11-54882.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[12]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_1[12]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_1[12]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54876.11-54882.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[12]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_2[12]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_2[12]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54883.11-54889.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[13]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_0[13]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_0[13]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54883.11-54889.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[13]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_1[13]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_1[13]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54883.11-54889.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[13]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_2[13]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_2[13]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54890.11-54896.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[14]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_0[14]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_0[14]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54890.11-54896.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[14]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_1[14]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_1[14]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54890.11-54896.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[14]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_2[14]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_2[14]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54897.11-54903.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[15]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_0[15]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_0[15]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54897.11-54903.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[15]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_1[15]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_1[15]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54897.11-54903.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[15]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_2[15]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_2[15]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54904.11-54910.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[16]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_0[16]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_0[16]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54904.11-54910.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[16]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_1[16]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_1[16]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54904.11-54910.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[16]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_2[16]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_2[16]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54911.11-54917.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[17]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_0[17]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_0[17]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54911.11-54917.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[17]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_1[17]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_1[17]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54911.11-54917.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[17]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_2[17]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_2[17]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54918.11-54924.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[18]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_0[18]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_0[18]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54918.11-54924.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[18]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_1[18]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_1[18]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54918.11-54924.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[18]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_2[18]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_2[18]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54925.11-54931.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[19]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_0[19]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_0[19]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54925.11-54931.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[19]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_1[19]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_1[19]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54925.11-54931.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[19]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_2[19]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_2[19]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54799.11-54805.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[1]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_0[1]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_0[1]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54799.11-54805.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[1]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_1[1]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_1[1]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54799.11-54805.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[1]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_2[1]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_2[1]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54932.11-54938.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[20]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_0[20]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_0[20]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54932.11-54938.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[20]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_1[20]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_1[20]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54932.11-54938.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[20]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_2[20]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_2[20]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54939.11-54945.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[21]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_0[21]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_0[21]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54939.11-54945.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[21]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_1[21]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_1[21]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54939.11-54945.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[21]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_2[21]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_2[21]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54946.11-54952.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[22]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_0[22]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_0[22]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54946.11-54952.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[22]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_1[22]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_1[22]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54946.11-54952.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[22]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_2[22]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_2[22]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54953.11-54959.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[23]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_0[23]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_0[23]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54953.11-54959.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[23]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_1[23]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_1[23]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54953.11-54959.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[23]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_2[23]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_2[23]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54960.11-54966.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[24]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_0[24]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_0[24]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54960.11-54966.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[24]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_1[24]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_1[24]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54960.11-54966.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[24]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_2[24]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_2[24]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54967.11-54973.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[25]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_0[25]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_0[25]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54967.11-54973.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[25]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_1[25]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_1[25]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54967.11-54973.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[25]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_2[25]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_2[25]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54974.11-54980.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[26]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_0[26]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_0[26]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54974.11-54980.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[26]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_1[26]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_1[26]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54974.11-54980.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[26]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_2[26]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_2[26]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54981.11-54987.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[27]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_0[27]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_0[27]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54981.11-54987.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[27]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_1[27]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_1[27]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54981.11-54987.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[27]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_2[27]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_2[27]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54988.11-54994.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[28]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_0[28]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_0[28]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54988.11-54994.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[28]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_1[28]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_1[28]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54988.11-54994.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[28]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_2[28]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_2[28]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54995.11-55001.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[29]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_0[29]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_0[29]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54995.11-55001.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[29]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_1[29]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_1[29]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54995.11-55001.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[29]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_2[29]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_2[29]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54806.11-54812.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[2]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_0[2]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_0[2]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54806.11-54812.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[2]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_1[2]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_1[2]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54806.11-54812.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[2]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_2[2]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_2[2]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55002.11-55008.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[30]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_0[30]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_0[30]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55002.11-55008.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[30]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_1[30]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_1[30]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55002.11-55008.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[30]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_2[30]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_2[30]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55009.11-55015.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[31]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_0[31]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_0[31]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55009.11-55015.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[31]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_1[31]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_1[31]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55009.11-55015.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[31]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_2[31]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_2[31]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54813.11-54819.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[3]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_0[3]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_0[3]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54813.11-54819.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[3]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_1[3]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_1[3]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54813.11-54819.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[3]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_2[3]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_2[3]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54820.11-54826.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[4]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_0[4]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_0[4]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54820.11-54826.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[4]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_1[4]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_1[4]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54820.11-54826.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[4]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_2[4]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_2[4]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54827.11-54833.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[5]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_0[5]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_0[5]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54827.11-54833.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[5]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_1[5]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_1[5]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54827.11-54833.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[5]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_2[5]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_2[5]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54834.11-54840.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[6]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_0[6]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_0[6]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54834.11-54840.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[6]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_1[6]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_1[6]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54834.11-54840.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[6]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_2[6]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_2[6]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54841.11-54847.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[7]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_0[7]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_0[7]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54841.11-54847.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[7]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_1[7]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_1[7]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54841.11-54847.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[7]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_2[7]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_2[7]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54848.11-54854.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[8]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_0[8]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_0[8]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54848.11-54854.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[8]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_1[8]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_1[8]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54848.11-54854.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[8]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_2[8]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_2[8]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54855.11-54861.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[9]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_0[9]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_0[9]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54855.11-54861.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[9]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_1[9]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_1[9]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54855.11-54861.2" *)
  FD1P3IX \builder_csr_bankarray_interface2_bank_bus_dat_r_reg[9]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface2_bank_bus_dat_r_11_TMR_2[9]),
    .Q(builder_csr_bankarray_interface2_bank_bus_dat_r_TMR_2[9]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54736.11-54742.2" *)
  FD1P3IX \builder_csr_bankarray_interface3_bank_bus_dat_r_reg[0]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface3_bank_bus_dat_r_11_TMR_0[0]),
    .Q(builder_csr_bankarray_interface3_bank_bus_dat_r_TMR_0[0]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54736.11-54742.2" *)
  FD1P3IX \builder_csr_bankarray_interface3_bank_bus_dat_r_reg[0]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface3_bank_bus_dat_r_11_TMR_1[0]),
    .Q(builder_csr_bankarray_interface3_bank_bus_dat_r_TMR_1[0]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54736.11-54742.2" *)
  FD1P3IX \builder_csr_bankarray_interface3_bank_bus_dat_r_reg[0]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface3_bank_bus_dat_r_11_TMR_2[0]),
    .Q(builder_csr_bankarray_interface3_bank_bus_dat_r_TMR_2[0]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54743.11-54749.2" *)
  FD1P3IX \builder_csr_bankarray_interface3_bank_bus_dat_r_reg[1]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface3_bank_bus_dat_r_11_TMR_0[1]),
    .Q(builder_csr_bankarray_interface3_bank_bus_dat_r_TMR_0[1]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54743.11-54749.2" *)
  FD1P3IX \builder_csr_bankarray_interface3_bank_bus_dat_r_reg[1]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface3_bank_bus_dat_r_11_TMR_1[1]),
    .Q(builder_csr_bankarray_interface3_bank_bus_dat_r_TMR_1[1]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54743.11-54749.2" *)
  FD1P3IX \builder_csr_bankarray_interface3_bank_bus_dat_r_reg[1]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_interface3_bank_bus_dat_r_11_TMR_2[1]),
    .Q(builder_csr_bankarray_interface3_bank_bus_dat_r_TMR_2[1]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54750.11-54756.2" *)
  FD1P3IX \builder_csr_bankarray_interface3_bank_bus_dat_r_reg[2]_TMR_0  (
    .CD(builder_csr_bankarray_interface3_bank_bus_dat_r_0_sqmuxa_i_TMR_0),
    .CK(sys_clk),
    .D(storage_1_dat1_TMR_0[2]),
    .Q(builder_csr_bankarray_interface3_bank_bus_dat_r_TMR_0[2]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54750.11-54756.2" *)
  FD1P3IX \builder_csr_bankarray_interface3_bank_bus_dat_r_reg[2]_TMR_1  (
    .CD(builder_csr_bankarray_interface3_bank_bus_dat_r_0_sqmuxa_i_TMR_1),
    .CK(sys_clk),
    .D(storage_1_dat1_TMR_1[2]),
    .Q(builder_csr_bankarray_interface3_bank_bus_dat_r_TMR_1[2]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54750.11-54756.2" *)
  FD1P3IX \builder_csr_bankarray_interface3_bank_bus_dat_r_reg[2]_TMR_2  (
    .CD(builder_csr_bankarray_interface3_bank_bus_dat_r_0_sqmuxa_i_TMR_2),
    .CK(sys_clk),
    .D(storage_1_dat1_TMR_2[2]),
    .Q(builder_csr_bankarray_interface3_bank_bus_dat_r_TMR_2[2]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54757.11-54763.2" *)
  FD1P3IX \builder_csr_bankarray_interface3_bank_bus_dat_r_reg[3]_TMR_0  (
    .CD(builder_csr_bankarray_interface3_bank_bus_dat_r_0_sqmuxa_i_TMR_0),
    .CK(sys_clk),
    .D(storage_1_dat1_TMR_0[3]),
    .Q(builder_csr_bankarray_interface3_bank_bus_dat_r_TMR_0[3]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54757.11-54763.2" *)
  FD1P3IX \builder_csr_bankarray_interface3_bank_bus_dat_r_reg[3]_TMR_1  (
    .CD(builder_csr_bankarray_interface3_bank_bus_dat_r_0_sqmuxa_i_TMR_1),
    .CK(sys_clk),
    .D(storage_1_dat1_TMR_1[3]),
    .Q(builder_csr_bankarray_interface3_bank_bus_dat_r_TMR_1[3]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54757.11-54763.2" *)
  FD1P3IX \builder_csr_bankarray_interface3_bank_bus_dat_r_reg[3]_TMR_2  (
    .CD(builder_csr_bankarray_interface3_bank_bus_dat_r_0_sqmuxa_i_TMR_2),
    .CK(sys_clk),
    .D(storage_1_dat1_TMR_2[3]),
    .Q(builder_csr_bankarray_interface3_bank_bus_dat_r_TMR_2[3]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54764.11-54770.2" *)
  FD1P3IX \builder_csr_bankarray_interface3_bank_bus_dat_r_reg[4]_TMR_0  (
    .CD(builder_csr_bankarray_interface3_bank_bus_dat_r_0_sqmuxa_i_TMR_0),
    .CK(sys_clk),
    .D(storage_1_dat1_TMR_0[4]),
    .Q(builder_csr_bankarray_interface3_bank_bus_dat_r_TMR_0[4]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54764.11-54770.2" *)
  FD1P3IX \builder_csr_bankarray_interface3_bank_bus_dat_r_reg[4]_TMR_1  (
    .CD(builder_csr_bankarray_interface3_bank_bus_dat_r_0_sqmuxa_i_TMR_1),
    .CK(sys_clk),
    .D(storage_1_dat1_TMR_1[4]),
    .Q(builder_csr_bankarray_interface3_bank_bus_dat_r_TMR_1[4]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54764.11-54770.2" *)
  FD1P3IX \builder_csr_bankarray_interface3_bank_bus_dat_r_reg[4]_TMR_2  (
    .CD(builder_csr_bankarray_interface3_bank_bus_dat_r_0_sqmuxa_i_TMR_2),
    .CK(sys_clk),
    .D(storage_1_dat1_TMR_2[4]),
    .Q(builder_csr_bankarray_interface3_bank_bus_dat_r_TMR_2[4]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54771.11-54777.2" *)
  FD1P3IX \builder_csr_bankarray_interface3_bank_bus_dat_r_reg[5]_TMR_0  (
    .CD(builder_csr_bankarray_interface3_bank_bus_dat_r_0_sqmuxa_i_TMR_0),
    .CK(sys_clk),
    .D(storage_1_dat1_TMR_0[5]),
    .Q(builder_csr_bankarray_interface3_bank_bus_dat_r_TMR_0[5]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54771.11-54777.2" *)
  FD1P3IX \builder_csr_bankarray_interface3_bank_bus_dat_r_reg[5]_TMR_1  (
    .CD(builder_csr_bankarray_interface3_bank_bus_dat_r_0_sqmuxa_i_TMR_1),
    .CK(sys_clk),
    .D(storage_1_dat1_TMR_1[5]),
    .Q(builder_csr_bankarray_interface3_bank_bus_dat_r_TMR_1[5]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54771.11-54777.2" *)
  FD1P3IX \builder_csr_bankarray_interface3_bank_bus_dat_r_reg[5]_TMR_2  (
    .CD(builder_csr_bankarray_interface3_bank_bus_dat_r_0_sqmuxa_i_TMR_2),
    .CK(sys_clk),
    .D(storage_1_dat1_TMR_2[5]),
    .Q(builder_csr_bankarray_interface3_bank_bus_dat_r_TMR_2[5]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54778.11-54784.2" *)
  FD1P3IX \builder_csr_bankarray_interface3_bank_bus_dat_r_reg[6]_TMR_0  (
    .CD(builder_csr_bankarray_interface3_bank_bus_dat_r_0_sqmuxa_i_TMR_0),
    .CK(sys_clk),
    .D(storage_1_dat1_TMR_0[6]),
    .Q(builder_csr_bankarray_interface3_bank_bus_dat_r_TMR_0[6]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54778.11-54784.2" *)
  FD1P3IX \builder_csr_bankarray_interface3_bank_bus_dat_r_reg[6]_TMR_1  (
    .CD(builder_csr_bankarray_interface3_bank_bus_dat_r_0_sqmuxa_i_TMR_1),
    .CK(sys_clk),
    .D(storage_1_dat1_TMR_1[6]),
    .Q(builder_csr_bankarray_interface3_bank_bus_dat_r_TMR_1[6]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54778.11-54784.2" *)
  FD1P3IX \builder_csr_bankarray_interface3_bank_bus_dat_r_reg[6]_TMR_2  (
    .CD(builder_csr_bankarray_interface3_bank_bus_dat_r_0_sqmuxa_i_TMR_2),
    .CK(sys_clk),
    .D(storage_1_dat1_TMR_2[6]),
    .Q(builder_csr_bankarray_interface3_bank_bus_dat_r_TMR_2[6]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54785.11-54791.2" *)
  FD1P3IX \builder_csr_bankarray_interface3_bank_bus_dat_r_reg[7]_TMR_0  (
    .CD(builder_csr_bankarray_interface3_bank_bus_dat_r_0_sqmuxa_i_TMR_0),
    .CK(sys_clk),
    .D(storage_1_dat1_TMR_0[7]),
    .Q(builder_csr_bankarray_interface3_bank_bus_dat_r_TMR_0[7]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54785.11-54791.2" *)
  FD1P3IX \builder_csr_bankarray_interface3_bank_bus_dat_r_reg[7]_TMR_1  (
    .CD(builder_csr_bankarray_interface3_bank_bus_dat_r_0_sqmuxa_i_TMR_1),
    .CK(sys_clk),
    .D(storage_1_dat1_TMR_1[7]),
    .Q(builder_csr_bankarray_interface3_bank_bus_dat_r_TMR_1[7]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54785.11-54791.2" *)
  FD1P3IX \builder_csr_bankarray_interface3_bank_bus_dat_r_reg[7]_TMR_2  (
    .CD(builder_csr_bankarray_interface3_bank_bus_dat_r_0_sqmuxa_i_TMR_2),
    .CK(sys_clk),
    .D(storage_1_dat1_TMR_2[7]),
    .Q(builder_csr_bankarray_interface3_bank_bus_dat_r_TMR_2[7]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54729.11-54735.2" *)
  FD1P3IX builder_csr_bankarray_sel_r_reg_TMR_0 (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(builder_csr_bankarray_sel_r_r_0_a2_TMR_0),
    .Q(builder_csr_bankarray_sel_r_TMR_0),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54729.11-54735.2" *)
  FD1P3IX builder_csr_bankarray_sel_r_reg_TMR_1 (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(builder_csr_bankarray_sel_r_r_0_a2_TMR_1),
    .Q(builder_csr_bankarray_sel_r_TMR_1),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54729.11-54735.2" *)
  FD1P3IX builder_csr_bankarray_sel_r_reg_TMR_2 (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(builder_csr_bankarray_sel_r_r_0_a2_TMR_2),
    .Q(builder_csr_bankarray_sel_r_TMR_2),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54715.11-54721.2" *)
  FD1P3IX builder_grant_fast_reg_TMR_0 (
    .CD(GND_0),
    .CK(sys_clk),
    .D(N_1210_i_fast_TMR_0),
    .Q(builder_grant_fast_TMR_0),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54715.11-54721.2" *)
  FD1P3IX builder_grant_fast_reg_TMR_1 (
    .CD(GND_0),
    .CK(sys_clk),
    .D(N_1210_i_fast_TMR_1),
    .Q(builder_grant_fast_TMR_1),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54715.11-54721.2" *)
  FD1P3IX builder_grant_fast_reg_TMR_2 (
    .CD(GND_0),
    .CK(sys_clk),
    .D(N_1210_i_fast_TMR_2),
    .Q(builder_grant_fast_TMR_2),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54722.11-54728.2" *)
  FD1P3IX builder_grant_reg_TMR_0 (
    .CD(GND_0),
    .CK(sys_clk),
    .D(N_1210_i_TMR_0),
    .Q(builder_grant_TMR_0),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54722.11-54728.2" *)
  FD1P3IX builder_grant_reg_TMR_1 (
    .CD(GND_0),
    .CK(sys_clk),
    .D(N_1210_i_TMR_1),
    .Q(builder_grant_TMR_1),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54722.11-54728.2" *)
  FD1P3IX builder_grant_reg_TMR_2 (
    .CD(GND_0),
    .CK(sys_clk),
    .D(N_1210_i_TMR_2),
    .Q(builder_grant_TMR_2),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54708.11-54714.2" *)
  FD1P3IX builder_grant_rep1_reg_TMR_0 (
    .CD(GND_0),
    .CK(sys_clk),
    .D(N_1210_i_rep1_TMR_0),
    .Q(builder_grant_rep1_TMR_0),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54708.11-54714.2" *)
  FD1P3IX builder_grant_rep1_reg_TMR_1 (
    .CD(GND_0),
    .CK(sys_clk),
    .D(N_1210_i_rep1_TMR_1),
    .Q(builder_grant_rep1_TMR_1),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54708.11-54714.2" *)
  FD1P3IX builder_grant_rep1_reg_TMR_2 (
    .CD(GND_0),
    .CK(sys_clk),
    .D(N_1210_i_rep1_TMR_2),
    .Q(builder_grant_rep1_TMR_2),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54701.11-54707.2" *)
  FD1P3IX builder_grant_rep2_reg_TMR_0 (
    .CD(GND_0),
    .CK(sys_clk),
    .D(N_1210_i_rep2_TMR_0),
    .Q(builder_grant_rep2_TMR_0),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54701.11-54707.2" *)
  FD1P3IX builder_grant_rep2_reg_TMR_1 (
    .CD(GND_0),
    .CK(sys_clk),
    .D(N_1210_i_rep2_TMR_1),
    .Q(builder_grant_rep2_TMR_1),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54701.11-54707.2" *)
  FD1P3IX builder_grant_rep2_reg_TMR_2 (
    .CD(GND_0),
    .CK(sys_clk),
    .D(N_1210_i_rep2_TMR_2),
    .Q(builder_grant_rep2_TMR_2),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51675.12-51681.2" *)
  IFD1P3IX builder_regs0_0io_TMR_0 (
    .CD(GND_0),
    .CK(sys_clk),
    .D(serial_rx_c),
    .Q(builder_regs0_TMR_0),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51675.12-51681.2" *)
  IFD1P3IX builder_regs0_0io_TMR_1 (
    .CD(GND_0),
    .CK(sys_clk),
    .D(serial_rx_c),
    .Q(builder_regs0_TMR_1),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51675.12-51681.2" *)
  IFD1P3IX builder_regs0_0io_TMR_2 (
    .CD(GND_0),
    .CK(sys_clk),
    .D(serial_rx_c),
    .Q(builder_regs0_TMR_2),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54694.11-54700.2" *)
  FD1P3IX builder_regs1_reg_TMR_0 (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_regs0_TMR_0),
    .Q(builder_regs1_TMR_0),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54694.11-54700.2" *)
  FD1P3IX builder_regs1_reg_TMR_1 (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_regs0_TMR_1),
    .Q(builder_regs1_TMR_1),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54694.11-54700.2" *)
  FD1P3IX builder_regs1_reg_TMR_2 (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_regs0_TMR_2),
    .Q(builder_regs1_TMR_2),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54673.11-54679.2" *)
  FD1P3IX \builder_slave_sel_r_reg[0]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(builder_slave_sel_2_TMR_0),
    .Q(builder_slave_sel_r_TMR_0[0]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54673.11-54679.2" *)
  FD1P3IX \builder_slave_sel_r_reg[0]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(builder_slave_sel_2_TMR_1),
    .Q(builder_slave_sel_r_TMR_1[0]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54673.11-54679.2" *)
  FD1P3IX \builder_slave_sel_r_reg[0]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(builder_slave_sel_2_TMR_2),
    .Q(builder_slave_sel_r_TMR_2[0]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54680.11-54686.2" *)
  FD1P3IX \builder_slave_sel_r_reg[1]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_slave_sel_r_r_0_a2_TMR_0),
    .Q(builder_slave_sel_r_TMR_0[1]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54680.11-54686.2" *)
  FD1P3IX \builder_slave_sel_r_reg[1]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_slave_sel_r_r_0_a2_TMR_1),
    .Q(builder_slave_sel_r_TMR_1[1]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54680.11-54686.2" *)
  FD1P3IX \builder_slave_sel_r_reg[1]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_slave_sel_r_r_0_a2_TMR_2),
    .Q(builder_slave_sel_r_TMR_2[1]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54687.11-54693.2" *)
  FD1P3IX \builder_slave_sel_r_reg[2]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(N_175_TMR_0),
    .Q(builder_slave_sel_r_TMR_0[2]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54687.11-54693.2" *)
  FD1P3IX \builder_slave_sel_r_reg[2]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(N_175_TMR_1),
    .Q(builder_slave_sel_r_TMR_1[2]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54687.11-54693.2" *)
  FD1P3IX \builder_slave_sel_r_reg[2]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(N_175_TMR_2),
    .Q(builder_slave_sel_r_TMR_2[2]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55573.6-55576.2" *)
  IB gsrn_pad (
    .I(gsrn),
    .O(gsrn_c)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51294.7-51297.2" *)
  INV gsrn_pad_RNIED4D_TMR_0 (
    .A(gsrn_c),
    .Z(gsrn_c_i_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51294.7-51297.2" *)
  INV gsrn_pad_RNIED4D_TMR_1 (
    .A(gsrn_c),
    .Z(gsrn_c_i_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51294.7-51297.2" *)
  INV gsrn_pad_RNIED4D_TMR_2 (
    .A(gsrn_c),
    .Z(gsrn_c_i_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54666.11-54672.2" *)
  FD1P3IX \main_basesoc_bus_errors_0_mod[0]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_bus_errors_0_mod_RNO_TMR_0),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_0[0]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54666.11-54672.2" *)
  FD1P3IX \main_basesoc_bus_errors_0_mod[0]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_bus_errors_0_mod_RNO_TMR_1),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_1[0]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54666.11-54672.2" *)
  FD1P3IX \main_basesoc_bus_errors_0_mod[0]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_bus_errors_0_mod_RNO_TMR_2),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_2[0]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56066.8-56072.2" *)
  LUT4 \main_basesoc_bus_errors_0_mod_RNO_cZ[0]_TMR_0  (
    .A(sys_rst_TMR_0),
    .B(un1_main_basesoc_bus_errors_1_TMR_0[0]),
    .C(GND_0),
    .D(GND_0),
    .Z(main_basesoc_bus_errors_0_mod_RNO_TMR_0)
  );
  defparam \main_basesoc_bus_errors_0_mod_RNO_cZ[0]_TMR_0 .INIT = "0x4444";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56066.8-56072.2" *)
  LUT4 \main_basesoc_bus_errors_0_mod_RNO_cZ[0]_TMR_1  (
    .A(sys_rst_TMR_1),
    .B(un1_main_basesoc_bus_errors_1_TMR_1[0]),
    .C(GND_0),
    .D(GND_0),
    .Z(main_basesoc_bus_errors_0_mod_RNO_TMR_1)
  );
  defparam \main_basesoc_bus_errors_0_mod_RNO_cZ[0]_TMR_1 .INIT = "0x4444";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56066.8-56072.2" *)
  LUT4 \main_basesoc_bus_errors_0_mod_RNO_cZ[0]_TMR_2  (
    .A(sys_rst_TMR_2),
    .B(un1_main_basesoc_bus_errors_1_TMR_2[0]),
    .C(GND_0),
    .D(GND_0),
    .Z(main_basesoc_bus_errors_0_mod_RNO_TMR_2)
  );
  defparam \main_basesoc_bus_errors_0_mod_RNO_cZ[0]_TMR_2 .INIT = "0x4444";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54512.11-54518.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[10]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_0[10]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_0[10]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54512.11-54518.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[10]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_1[10]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_1[10]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54512.11-54518.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[10]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_2[10]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_2[10]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54519.11-54525.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[11]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_0[11]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_0[11]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54519.11-54525.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[11]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_1[11]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_1[11]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54519.11-54525.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[11]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_2[11]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_2[11]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54526.11-54532.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[12]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_0[12]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_0[12]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54526.11-54532.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[12]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_1[12]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_1[12]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54526.11-54532.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[12]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_2[12]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_2[12]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54533.11-54539.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[13]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_0[13]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_0[13]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54533.11-54539.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[13]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_1[13]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_1[13]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54533.11-54539.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[13]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_2[13]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_2[13]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54540.11-54546.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[14]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_0[14]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_0[14]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54540.11-54546.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[14]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_1[14]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_1[14]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54540.11-54546.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[14]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_2[14]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_2[14]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54547.11-54553.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[15]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_0[15]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_0[15]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54547.11-54553.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[15]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_1[15]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_1[15]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54547.11-54553.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[15]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_2[15]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_2[15]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54554.11-54560.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[16]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_0[16]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_0[16]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54554.11-54560.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[16]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_1[16]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_1[16]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54554.11-54560.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[16]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_2[16]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_2[16]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54561.11-54567.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[17]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_0[17]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_0[17]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54561.11-54567.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[17]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_1[17]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_1[17]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54561.11-54567.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[17]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_2[17]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_2[17]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54568.11-54574.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[18]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_0[18]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_0[18]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54568.11-54574.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[18]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_1[18]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_1[18]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54568.11-54574.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[18]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_2[18]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_2[18]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54575.11-54581.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[19]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_0[19]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_0[19]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54575.11-54581.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[19]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_1[19]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_1[19]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54575.11-54581.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[19]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_2[19]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_2[19]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54449.11-54455.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[1]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_0[1]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_0[1]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54449.11-54455.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[1]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_1[1]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_1[1]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54449.11-54455.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[1]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_2[1]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_2[1]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54582.11-54588.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[20]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_0[20]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_0[20]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54582.11-54588.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[20]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_1[20]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_1[20]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54582.11-54588.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[20]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_2[20]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_2[20]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54589.11-54595.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[21]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_0[21]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_0[21]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54589.11-54595.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[21]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_1[21]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_1[21]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54589.11-54595.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[21]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_2[21]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_2[21]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54596.11-54602.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[22]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_0[22]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_0[22]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54596.11-54602.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[22]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_1[22]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_1[22]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54596.11-54602.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[22]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_2[22]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_2[22]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54603.11-54609.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[23]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_0[23]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_0[23]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54603.11-54609.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[23]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_1[23]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_1[23]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54603.11-54609.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[23]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_2[23]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_2[23]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54610.11-54616.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[24]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_0[24]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_0[24]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54610.11-54616.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[24]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_1[24]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_1[24]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54610.11-54616.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[24]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_2[24]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_2[24]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54617.11-54623.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[25]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_0[25]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_0[25]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54617.11-54623.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[25]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_1[25]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_1[25]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54617.11-54623.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[25]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_2[25]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_2[25]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54624.11-54630.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[26]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_0[26]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_0[26]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54624.11-54630.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[26]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_1[26]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_1[26]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54624.11-54630.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[26]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_2[26]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_2[26]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54631.11-54637.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[27]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_0[27]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_0[27]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54631.11-54637.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[27]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_1[27]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_1[27]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54631.11-54637.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[27]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_2[27]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_2[27]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54638.11-54644.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[28]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_0[28]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_0[28]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54638.11-54644.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[28]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_1[28]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_1[28]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54638.11-54644.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[28]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_2[28]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_2[28]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54645.11-54651.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[29]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_0[29]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_0[29]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54645.11-54651.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[29]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_1[29]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_1[29]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54645.11-54651.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[29]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_2[29]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_2[29]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54456.11-54462.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[2]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_0[2]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_0[2]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54456.11-54462.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[2]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_1[2]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_1[2]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54456.11-54462.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[2]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_2[2]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_2[2]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54652.11-54658.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[30]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_0[30]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_0[30]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54652.11-54658.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[30]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_1[30]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_1[30]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54652.11-54658.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[30]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_2[30]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_2[30]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54659.11-54665.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[31]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_0[31]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_0[31]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54659.11-54665.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[31]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_1[31]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_1[31]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54659.11-54665.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[31]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_2[31]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_2[31]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54463.11-54469.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[3]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_0[3]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_0[3]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54463.11-54469.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[3]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_1[3]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_1[3]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54463.11-54469.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[3]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_2[3]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_2[3]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54470.11-54476.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[4]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_0[4]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_0[4]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54470.11-54476.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[4]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_1[4]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_1[4]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54470.11-54476.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[4]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_2[4]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_2[4]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54477.11-54483.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[5]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_0[5]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_0[5]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54477.11-54483.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[5]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_1[5]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_1[5]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54477.11-54483.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[5]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_2[5]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_2[5]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54484.11-54490.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[6]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_0[6]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_0[6]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54484.11-54490.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[6]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_1[6]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_1[6]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54484.11-54490.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[6]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_2[6]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_2[6]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54491.11-54497.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[7]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_0[7]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_0[7]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54491.11-54497.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[7]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_1[7]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_1[7]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54491.11-54497.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[7]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_2[7]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_2[7]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54498.11-54504.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[8]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_0[8]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_0[8]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54498.11-54504.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[8]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_1[8]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_1[8]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54498.11-54504.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[8]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_2[8]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_2[8]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54505.11-54511.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[9]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_0[9]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_0[9]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54505.11-54511.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[9]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_1[9]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_1[9]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54505.11-54511.2" *)
  FD1P3IX \main_basesoc_bus_errors_mod[9]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_bus_errors_1_TMR_2[9]),
    .Q(un1_main_basesoc_bus_errors_1_0_TMR_2[9]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54442.11-54448.2" *)
  FD1P3IX main_basesoc_ram_bus_ack_reg_TMR_0 (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(main_basesoc_ram_bus_ack_r_TMR_0),
    .Q(main_basesoc_ram_bus_ack_TMR_0),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54442.11-54448.2" *)
  FD1P3IX main_basesoc_ram_bus_ack_reg_TMR_1 (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(main_basesoc_ram_bus_ack_r_TMR_1),
    .Q(main_basesoc_ram_bus_ack_TMR_1),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54442.11-54448.2" *)
  FD1P3IX main_basesoc_ram_bus_ack_reg_TMR_2 (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(main_basesoc_ram_bus_ack_r_TMR_2),
    .Q(main_basesoc_ram_bus_ack_TMR_2),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54435.11-54441.2" *)
  FD1P3IX main_basesoc_reset_re_reg_TMR_0 (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_reset_storage_0_sqmuxa_TMR_0),
    .Q(main_basesoc_reset_re_TMR_0),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54435.11-54441.2" *)
  FD1P3IX main_basesoc_reset_re_reg_TMR_1 (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_reset_storage_0_sqmuxa_TMR_1),
    .Q(main_basesoc_reset_re_TMR_1),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54435.11-54441.2" *)
  FD1P3IX main_basesoc_reset_re_reg_TMR_2 (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_reset_storage_0_sqmuxa_TMR_2),
    .Q(main_basesoc_reset_re_TMR_2),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54421.11-54427.2" *)
  FD1P3IX \main_basesoc_reset_storage_reg[0]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[0]),
    .Q(main_basesoc_reset_storage_TMR_0[0]),
    .SP(builder_csr_bankarray_csrbank0_reset0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54421.11-54427.2" *)
  FD1P3IX \main_basesoc_reset_storage_reg[0]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[0]),
    .Q(main_basesoc_reset_storage_TMR_1[0]),
    .SP(builder_csr_bankarray_csrbank0_reset0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54421.11-54427.2" *)
  FD1P3IX \main_basesoc_reset_storage_reg[0]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[0]),
    .Q(main_basesoc_reset_storage_TMR_2[0]),
    .SP(builder_csr_bankarray_csrbank0_reset0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54428.11-54434.2" *)
  FD1P3IX \main_basesoc_reset_storage_reg[1]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[1]),
    .Q(main_basesoc_reset_storage_TMR_0[1]),
    .SP(builder_csr_bankarray_csrbank0_reset0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54428.11-54434.2" *)
  FD1P3IX \main_basesoc_reset_storage_reg[1]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[1]),
    .Q(main_basesoc_reset_storage_TMR_1[1]),
    .SP(builder_csr_bankarray_csrbank0_reset0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54428.11-54434.2" *)
  FD1P3IX \main_basesoc_reset_storage_reg[1]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[1]),
    .Q(main_basesoc_reset_storage_TMR_2[1]),
    .SP(builder_csr_bankarray_csrbank0_reset0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54393.11-54399.2" *)
  FD1P3IX \main_basesoc_rx_count[0]_TMR_0  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_0),
    .CK(sys_clk),
    .D(\main_basesoc_rx_count_0_.fb_TMR_0 ),
    .Q(CO0_TMR_0),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54393.11-54399.2" *)
  FD1P3IX \main_basesoc_rx_count[0]_TMR_1  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_1),
    .CK(sys_clk),
    .D(\main_basesoc_rx_count_0_.fb_TMR_1 ),
    .Q(CO0_TMR_1),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54393.11-54399.2" *)
  FD1P3IX \main_basesoc_rx_count[0]_TMR_2  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_2),
    .CK(sys_clk),
    .D(\main_basesoc_rx_count_0_.fb_TMR_2 ),
    .Q(CO0_TMR_2),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51389.8-51395.2" *)
  LUT4 \main_basesoc_rx_count_0_.fb_cZ_TMR_0  (
    .A(CO0_TMR_0),
    .B(main_basesoc_rx_tick_TMR_0),
    .C(builder_basesoc_rs232phyrx_state_TMR_0),
    .D(GND_0),
    .Z(\main_basesoc_rx_count_0_.fb_TMR_0 )
  );
  defparam \main_basesoc_rx_count_0_.fb_cZ_TMR_0 .INIT = "0x6565";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51389.8-51395.2" *)
  LUT4 \main_basesoc_rx_count_0_.fb_cZ_TMR_1  (
    .A(CO0_TMR_1),
    .B(main_basesoc_rx_tick_TMR_1),
    .C(builder_basesoc_rs232phyrx_state_TMR_1),
    .D(GND_0),
    .Z(\main_basesoc_rx_count_0_.fb_TMR_1 )
  );
  defparam \main_basesoc_rx_count_0_.fb_cZ_TMR_1 .INIT = "0x6565";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51389.8-51395.2" *)
  LUT4 \main_basesoc_rx_count_0_.fb_cZ_TMR_2  (
    .A(CO0_TMR_2),
    .B(main_basesoc_rx_tick_TMR_2),
    .C(builder_basesoc_rs232phyrx_state_TMR_2),
    .D(GND_0),
    .Z(\main_basesoc_rx_count_0_.fb_TMR_2 )
  );
  defparam \main_basesoc_rx_count_0_.fb_cZ_TMR_2 .INIT = "0x6565";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54400.11-54406.2" *)
  FD1P3IX \main_basesoc_rx_count_reg[1]_TMR_0  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_0),
    .CK(sys_clk),
    .D(main_basesoc_rx_count_rs232phyrx_next_value0_TMR_0[1]),
    .Q(main_basesoc_rx_count_TMR_0[1]),
    .SP(main_basesoc_rx_count_rs232phyrx_next_value_ce0_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54400.11-54406.2" *)
  FD1P3IX \main_basesoc_rx_count_reg[1]_TMR_1  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_1),
    .CK(sys_clk),
    .D(main_basesoc_rx_count_rs232phyrx_next_value0_TMR_1[1]),
    .Q(main_basesoc_rx_count_TMR_1[1]),
    .SP(main_basesoc_rx_count_rs232phyrx_next_value_ce0_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54400.11-54406.2" *)
  FD1P3IX \main_basesoc_rx_count_reg[1]_TMR_2  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_2),
    .CK(sys_clk),
    .D(main_basesoc_rx_count_rs232phyrx_next_value0_TMR_2[1]),
    .Q(main_basesoc_rx_count_TMR_2[1]),
    .SP(main_basesoc_rx_count_rs232phyrx_next_value_ce0_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54407.11-54413.2" *)
  FD1P3IX \main_basesoc_rx_count_reg[2]_TMR_0  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_0),
    .CK(sys_clk),
    .D(main_basesoc_rx_count_rs232phyrx_next_value0_TMR_0[2]),
    .Q(main_basesoc_rx_count_TMR_0[2]),
    .SP(main_basesoc_rx_count_rs232phyrx_next_value_ce0_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54407.11-54413.2" *)
  FD1P3IX \main_basesoc_rx_count_reg[2]_TMR_1  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_1),
    .CK(sys_clk),
    .D(main_basesoc_rx_count_rs232phyrx_next_value0_TMR_1[2]),
    .Q(main_basesoc_rx_count_TMR_1[2]),
    .SP(main_basesoc_rx_count_rs232phyrx_next_value_ce0_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54407.11-54413.2" *)
  FD1P3IX \main_basesoc_rx_count_reg[2]_TMR_2  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_2),
    .CK(sys_clk),
    .D(main_basesoc_rx_count_rs232phyrx_next_value0_TMR_2[2]),
    .Q(main_basesoc_rx_count_TMR_2[2]),
    .SP(main_basesoc_rx_count_rs232phyrx_next_value_ce0_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54414.11-54420.2" *)
  FD1P3IX \main_basesoc_rx_count_reg[3]_TMR_0  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_0),
    .CK(sys_clk),
    .D(main_basesoc_rx_count_rs232phyrx_next_value0_TMR_0[3]),
    .Q(main_basesoc_rx_count_TMR_0[3]),
    .SP(main_basesoc_rx_count_rs232phyrx_next_value_ce0_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54414.11-54420.2" *)
  FD1P3IX \main_basesoc_rx_count_reg[3]_TMR_1  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_1),
    .CK(sys_clk),
    .D(main_basesoc_rx_count_rs232phyrx_next_value0_TMR_1[3]),
    .Q(main_basesoc_rx_count_TMR_1[3]),
    .SP(main_basesoc_rx_count_rs232phyrx_next_value_ce0_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54414.11-54420.2" *)
  FD1P3IX \main_basesoc_rx_count_reg[3]_TMR_2  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_2),
    .CK(sys_clk),
    .D(main_basesoc_rx_count_rs232phyrx_next_value0_TMR_2[3]),
    .Q(main_basesoc_rx_count_TMR_2[3]),
    .SP(main_basesoc_rx_count_rs232phyrx_next_value_ce0_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54337.11-54343.2" *)
  FD1P3IX \main_basesoc_rx_data_reg[0]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_rx_data_TMR_0[1]),
    .Q(main_basesoc_rx_data_TMR_0[0]),
    .SP(main_basesoc_rx_data_rs232phyrx_next_value1_0_sqmuxa_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54337.11-54343.2" *)
  FD1P3IX \main_basesoc_rx_data_reg[0]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_rx_data_TMR_1[1]),
    .Q(main_basesoc_rx_data_TMR_1[0]),
    .SP(main_basesoc_rx_data_rs232phyrx_next_value1_0_sqmuxa_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54337.11-54343.2" *)
  FD1P3IX \main_basesoc_rx_data_reg[0]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_rx_data_TMR_2[1]),
    .Q(main_basesoc_rx_data_TMR_2[0]),
    .SP(main_basesoc_rx_data_rs232phyrx_next_value1_0_sqmuxa_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54344.11-54350.2" *)
  FD1P3IX \main_basesoc_rx_data_reg[1]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_rx_data_TMR_0[2]),
    .Q(main_basesoc_rx_data_TMR_0[1]),
    .SP(main_basesoc_rx_data_rs232phyrx_next_value1_0_sqmuxa_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54344.11-54350.2" *)
  FD1P3IX \main_basesoc_rx_data_reg[1]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_rx_data_TMR_1[2]),
    .Q(main_basesoc_rx_data_TMR_1[1]),
    .SP(main_basesoc_rx_data_rs232phyrx_next_value1_0_sqmuxa_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54344.11-54350.2" *)
  FD1P3IX \main_basesoc_rx_data_reg[1]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_rx_data_TMR_2[2]),
    .Q(main_basesoc_rx_data_TMR_2[1]),
    .SP(main_basesoc_rx_data_rs232phyrx_next_value1_0_sqmuxa_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54351.11-54357.2" *)
  FD1P3IX \main_basesoc_rx_data_reg[2]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_rx_data_TMR_0[3]),
    .Q(main_basesoc_rx_data_TMR_0[2]),
    .SP(main_basesoc_rx_data_rs232phyrx_next_value1_0_sqmuxa_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54351.11-54357.2" *)
  FD1P3IX \main_basesoc_rx_data_reg[2]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_rx_data_TMR_1[3]),
    .Q(main_basesoc_rx_data_TMR_1[2]),
    .SP(main_basesoc_rx_data_rs232phyrx_next_value1_0_sqmuxa_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54351.11-54357.2" *)
  FD1P3IX \main_basesoc_rx_data_reg[2]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_rx_data_TMR_2[3]),
    .Q(main_basesoc_rx_data_TMR_2[2]),
    .SP(main_basesoc_rx_data_rs232phyrx_next_value1_0_sqmuxa_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54358.11-54364.2" *)
  FD1P3IX \main_basesoc_rx_data_reg[3]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_rx_data_TMR_0[4]),
    .Q(main_basesoc_rx_data_TMR_0[3]),
    .SP(main_basesoc_rx_data_rs232phyrx_next_value1_0_sqmuxa_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54358.11-54364.2" *)
  FD1P3IX \main_basesoc_rx_data_reg[3]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_rx_data_TMR_1[4]),
    .Q(main_basesoc_rx_data_TMR_1[3]),
    .SP(main_basesoc_rx_data_rs232phyrx_next_value1_0_sqmuxa_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54358.11-54364.2" *)
  FD1P3IX \main_basesoc_rx_data_reg[3]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_rx_data_TMR_2[4]),
    .Q(main_basesoc_rx_data_TMR_2[3]),
    .SP(main_basesoc_rx_data_rs232phyrx_next_value1_0_sqmuxa_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54365.11-54371.2" *)
  FD1P3IX \main_basesoc_rx_data_reg[4]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_rx_data_TMR_0[5]),
    .Q(main_basesoc_rx_data_TMR_0[4]),
    .SP(main_basesoc_rx_data_rs232phyrx_next_value1_0_sqmuxa_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54365.11-54371.2" *)
  FD1P3IX \main_basesoc_rx_data_reg[4]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_rx_data_TMR_1[5]),
    .Q(main_basesoc_rx_data_TMR_1[4]),
    .SP(main_basesoc_rx_data_rs232phyrx_next_value1_0_sqmuxa_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54365.11-54371.2" *)
  FD1P3IX \main_basesoc_rx_data_reg[4]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_rx_data_TMR_2[5]),
    .Q(main_basesoc_rx_data_TMR_2[4]),
    .SP(main_basesoc_rx_data_rs232phyrx_next_value1_0_sqmuxa_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54372.11-54378.2" *)
  FD1P3IX \main_basesoc_rx_data_reg[5]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_rx_data_TMR_0[6]),
    .Q(main_basesoc_rx_data_TMR_0[5]),
    .SP(main_basesoc_rx_data_rs232phyrx_next_value1_0_sqmuxa_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54372.11-54378.2" *)
  FD1P3IX \main_basesoc_rx_data_reg[5]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_rx_data_TMR_1[6]),
    .Q(main_basesoc_rx_data_TMR_1[5]),
    .SP(main_basesoc_rx_data_rs232phyrx_next_value1_0_sqmuxa_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54372.11-54378.2" *)
  FD1P3IX \main_basesoc_rx_data_reg[5]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_rx_data_TMR_2[6]),
    .Q(main_basesoc_rx_data_TMR_2[5]),
    .SP(main_basesoc_rx_data_rs232phyrx_next_value1_0_sqmuxa_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54379.11-54385.2" *)
  FD1P3IX \main_basesoc_rx_data_reg[6]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_rx_data_TMR_0[7]),
    .Q(main_basesoc_rx_data_TMR_0[6]),
    .SP(main_basesoc_rx_data_rs232phyrx_next_value1_0_sqmuxa_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54379.11-54385.2" *)
  FD1P3IX \main_basesoc_rx_data_reg[6]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_rx_data_TMR_1[7]),
    .Q(main_basesoc_rx_data_TMR_1[6]),
    .SP(main_basesoc_rx_data_rs232phyrx_next_value1_0_sqmuxa_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54379.11-54385.2" *)
  FD1P3IX \main_basesoc_rx_data_reg[6]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_rx_data_TMR_2[7]),
    .Q(main_basesoc_rx_data_TMR_2[6]),
    .SP(main_basesoc_rx_data_rs232phyrx_next_value1_0_sqmuxa_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54386.11-54392.2" *)
  FD1P3IX \main_basesoc_rx_data_reg[7]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_regs1_TMR_0),
    .Q(main_basesoc_rx_data_TMR_0[7]),
    .SP(main_basesoc_rx_data_rs232phyrx_next_value1_0_sqmuxa_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54386.11-54392.2" *)
  FD1P3IX \main_basesoc_rx_data_reg[7]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_regs1_TMR_1),
    .Q(main_basesoc_rx_data_TMR_1[7]),
    .SP(main_basesoc_rx_data_rs232phyrx_next_value1_0_sqmuxa_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54386.11-54392.2" *)
  FD1P3IX \main_basesoc_rx_data_reg[7]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(builder_regs1_TMR_2),
    .Q(main_basesoc_rx_data_TMR_2[7]),
    .SP(main_basesoc_rx_data_rs232phyrx_next_value1_0_sqmuxa_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54330.11-54336.2" *)
  FD1P3IX \main_basesoc_rx_phase[31]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(N_17837_0_TMR_0),
    .Q(dsp_join_kb_27_TMR_0[31]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54330.11-54336.2" *)
  FD1P3IX \main_basesoc_rx_phase[31]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(N_17837_0_TMR_1),
    .Q(dsp_join_kb_27_TMR_1[31]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54330.11-54336.2" *)
  FD1P3IX \main_basesoc_rx_phase[31]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(N_17837_0_TMR_2),
    .Q(dsp_join_kb_27_TMR_2[31]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51667.8-51673.2" *)
  LUT4 \main_basesoc_rx_phase_RNO[31]_TMR_0  (
    .A(builder_basesoc_rs232phyrx_state_TMR_0),
    .B(un5_main_basesoc_rx_phase_cry_31_0_S0_TMR_0),
    .C(GND_0),
    .D(GND_0),
    .Z(N_17837_0_TMR_0)
  );
  defparam \main_basesoc_rx_phase_RNO[31]_TMR_0 .INIT = "0xDDDD";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51667.8-51673.2" *)
  LUT4 \main_basesoc_rx_phase_RNO[31]_TMR_1  (
    .A(builder_basesoc_rs232phyrx_state_TMR_1),
    .B(un5_main_basesoc_rx_phase_cry_31_0_S0_TMR_1),
    .C(GND_0),
    .D(GND_0),
    .Z(N_17837_0_TMR_1)
  );
  defparam \main_basesoc_rx_phase_RNO[31]_TMR_1 .INIT = "0xDDDD";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51667.8-51673.2" *)
  LUT4 \main_basesoc_rx_phase_RNO[31]_TMR_2  (
    .A(builder_basesoc_rs232phyrx_state_TMR_2),
    .B(un5_main_basesoc_rx_phase_cry_31_0_S0_TMR_2),
    .C(GND_0),
    .D(GND_0),
    .Z(N_17837_0_TMR_2)
  );
  defparam \main_basesoc_rx_phase_RNO[31]_TMR_2 .INIT = "0xDDDD";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54113.11-54119.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[0]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_rx_phase_mod_RNO_TMR_0),
    .Q(dsp_join_kb_27_TMR_0[0]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54113.11-54119.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[0]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_rx_phase_mod_RNO_TMR_1),
    .Q(dsp_join_kb_27_TMR_1[0]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54113.11-54119.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[0]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_rx_phase_mod_RNO_TMR_2),
    .Q(dsp_join_kb_27_TMR_2[0]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54183.11-54189.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[10]_TMR_0  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_0),
    .CK(sys_clk),
    .D(N_412_TMR_0),
    .Q(dsp_join_kb_27_TMR_0[10]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54183.11-54189.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[10]_TMR_1  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_1),
    .CK(sys_clk),
    .D(N_412_TMR_1),
    .Q(dsp_join_kb_27_TMR_1[10]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54183.11-54189.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[10]_TMR_2  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_2),
    .CK(sys_clk),
    .D(N_412_TMR_2),
    .Q(dsp_join_kb_27_TMR_2[10]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54190.11-54196.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[11]_TMR_0  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_0),
    .CK(sys_clk),
    .D(N_413_TMR_0),
    .Q(dsp_join_kb_27_TMR_0[11]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54190.11-54196.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[11]_TMR_1  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_1),
    .CK(sys_clk),
    .D(N_413_TMR_1),
    .Q(dsp_join_kb_27_TMR_1[11]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54190.11-54196.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[11]_TMR_2  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_2),
    .CK(sys_clk),
    .D(N_413_TMR_2),
    .Q(dsp_join_kb_27_TMR_2[11]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54197.11-54203.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[12]_TMR_0  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_0),
    .CK(sys_clk),
    .D(N_414_TMR_0),
    .Q(dsp_join_kb_27_TMR_0[12]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54197.11-54203.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[12]_TMR_1  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_1),
    .CK(sys_clk),
    .D(N_414_TMR_1),
    .Q(dsp_join_kb_27_TMR_1[12]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54197.11-54203.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[12]_TMR_2  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_2),
    .CK(sys_clk),
    .D(N_414_TMR_2),
    .Q(dsp_join_kb_27_TMR_2[12]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54204.11-54210.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[13]_TMR_0  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_0),
    .CK(sys_clk),
    .D(N_415_TMR_0),
    .Q(dsp_join_kb_27_TMR_0[13]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54204.11-54210.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[13]_TMR_1  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_1),
    .CK(sys_clk),
    .D(N_415_TMR_1),
    .Q(dsp_join_kb_27_TMR_1[13]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54204.11-54210.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[13]_TMR_2  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_2),
    .CK(sys_clk),
    .D(N_415_TMR_2),
    .Q(dsp_join_kb_27_TMR_2[13]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54211.11-54217.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[14]_TMR_0  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_0),
    .CK(sys_clk),
    .D(N_416_TMR_0),
    .Q(dsp_join_kb_27_TMR_0[14]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54211.11-54217.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[14]_TMR_1  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_1),
    .CK(sys_clk),
    .D(N_416_TMR_1),
    .Q(dsp_join_kb_27_TMR_1[14]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54211.11-54217.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[14]_TMR_2  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_2),
    .CK(sys_clk),
    .D(N_416_TMR_2),
    .Q(dsp_join_kb_27_TMR_2[14]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54218.11-54224.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[15]_TMR_0  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_0),
    .CK(sys_clk),
    .D(N_417_TMR_0),
    .Q(dsp_join_kb_27_TMR_0[15]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54218.11-54224.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[15]_TMR_1  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_1),
    .CK(sys_clk),
    .D(N_417_TMR_1),
    .Q(dsp_join_kb_27_TMR_1[15]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54218.11-54224.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[15]_TMR_2  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_2),
    .CK(sys_clk),
    .D(N_417_TMR_2),
    .Q(dsp_join_kb_27_TMR_2[15]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54225.11-54231.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[16]_TMR_0  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_0),
    .CK(sys_clk),
    .D(un5_main_basesoc_rx_phase_cry_15_0_S1_TMR_0),
    .Q(dsp_join_kb_27_TMR_0[16]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54225.11-54231.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[16]_TMR_1  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_1),
    .CK(sys_clk),
    .D(un5_main_basesoc_rx_phase_cry_15_0_S1_TMR_1),
    .Q(dsp_join_kb_27_TMR_1[16]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54225.11-54231.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[16]_TMR_2  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_2),
    .CK(sys_clk),
    .D(un5_main_basesoc_rx_phase_cry_15_0_S1_TMR_2),
    .Q(dsp_join_kb_27_TMR_2[16]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54232.11-54238.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[17]_TMR_0  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_0),
    .CK(sys_clk),
    .D(N_419_TMR_0),
    .Q(dsp_join_kb_27_TMR_0[17]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54232.11-54238.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[17]_TMR_1  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_1),
    .CK(sys_clk),
    .D(N_419_TMR_1),
    .Q(dsp_join_kb_27_TMR_1[17]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54232.11-54238.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[17]_TMR_2  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_2),
    .CK(sys_clk),
    .D(N_419_TMR_2),
    .Q(dsp_join_kb_27_TMR_2[17]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54239.11-54245.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[18]_TMR_0  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_0),
    .CK(sys_clk),
    .D(N_420_TMR_0),
    .Q(dsp_join_kb_27_TMR_0[18]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54239.11-54245.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[18]_TMR_1  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_1),
    .CK(sys_clk),
    .D(N_420_TMR_1),
    .Q(dsp_join_kb_27_TMR_1[18]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54239.11-54245.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[18]_TMR_2  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_2),
    .CK(sys_clk),
    .D(N_420_TMR_2),
    .Q(dsp_join_kb_27_TMR_2[18]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54246.11-54252.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[19]_TMR_0  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_0),
    .CK(sys_clk),
    .D(un5_main_basesoc_rx_phase_cry_19_0_S0_TMR_0),
    .Q(dsp_join_kb_27_TMR_0[19]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54246.11-54252.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[19]_TMR_1  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_1),
    .CK(sys_clk),
    .D(un5_main_basesoc_rx_phase_cry_19_0_S0_TMR_1),
    .Q(dsp_join_kb_27_TMR_1[19]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54246.11-54252.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[19]_TMR_2  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_2),
    .CK(sys_clk),
    .D(un5_main_basesoc_rx_phase_cry_19_0_S0_TMR_2),
    .Q(dsp_join_kb_27_TMR_2[19]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54120.11-54126.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[1]_TMR_0  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_0),
    .CK(sys_clk),
    .D(N_403_TMR_0),
    .Q(dsp_join_kb_27_TMR_0[1]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54120.11-54126.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[1]_TMR_1  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_1),
    .CK(sys_clk),
    .D(N_403_TMR_1),
    .Q(dsp_join_kb_27_TMR_1[1]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54120.11-54126.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[1]_TMR_2  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_2),
    .CK(sys_clk),
    .D(N_403_TMR_2),
    .Q(dsp_join_kb_27_TMR_2[1]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54253.11-54259.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[20]_TMR_0  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_0),
    .CK(sys_clk),
    .D(un5_main_basesoc_rx_phase_cry_19_0_S1_TMR_0),
    .Q(dsp_join_kb_27_TMR_0[20]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54253.11-54259.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[20]_TMR_1  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_1),
    .CK(sys_clk),
    .D(un5_main_basesoc_rx_phase_cry_19_0_S1_TMR_1),
    .Q(dsp_join_kb_27_TMR_1[20]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54253.11-54259.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[20]_TMR_2  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_2),
    .CK(sys_clk),
    .D(un5_main_basesoc_rx_phase_cry_19_0_S1_TMR_2),
    .Q(dsp_join_kb_27_TMR_2[20]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54260.11-54266.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[21]_TMR_0  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_0),
    .CK(sys_clk),
    .D(N_423_TMR_0),
    .Q(dsp_join_kb_27_TMR_0[21]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54260.11-54266.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[21]_TMR_1  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_1),
    .CK(sys_clk),
    .D(N_423_TMR_1),
    .Q(dsp_join_kb_27_TMR_1[21]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54260.11-54266.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[21]_TMR_2  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_2),
    .CK(sys_clk),
    .D(N_423_TMR_2),
    .Q(dsp_join_kb_27_TMR_2[21]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54267.11-54273.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[22]_TMR_0  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_0),
    .CK(sys_clk),
    .D(N_424_TMR_0),
    .Q(dsp_join_kb_27_TMR_0[22]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54267.11-54273.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[22]_TMR_1  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_1),
    .CK(sys_clk),
    .D(N_424_TMR_1),
    .Q(dsp_join_kb_27_TMR_1[22]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54267.11-54273.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[22]_TMR_2  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_2),
    .CK(sys_clk),
    .D(N_424_TMR_2),
    .Q(dsp_join_kb_27_TMR_2[22]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54274.11-54280.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[23]_TMR_0  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_0),
    .CK(sys_clk),
    .D(N_425_TMR_0),
    .Q(dsp_join_kb_27_TMR_0[23]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54274.11-54280.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[23]_TMR_1  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_1),
    .CK(sys_clk),
    .D(N_425_TMR_1),
    .Q(dsp_join_kb_27_TMR_1[23]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54274.11-54280.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[23]_TMR_2  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_2),
    .CK(sys_clk),
    .D(N_425_TMR_2),
    .Q(dsp_join_kb_27_TMR_2[23]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54281.11-54287.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[24]_TMR_0  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_0),
    .CK(sys_clk),
    .D(un5_main_basesoc_rx_phase_cry_23_0_S1_TMR_0),
    .Q(dsp_join_kb_27_TMR_0[24]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54281.11-54287.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[24]_TMR_1  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_1),
    .CK(sys_clk),
    .D(un5_main_basesoc_rx_phase_cry_23_0_S1_TMR_1),
    .Q(dsp_join_kb_27_TMR_1[24]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54281.11-54287.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[24]_TMR_2  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_2),
    .CK(sys_clk),
    .D(un5_main_basesoc_rx_phase_cry_23_0_S1_TMR_2),
    .Q(dsp_join_kb_27_TMR_2[24]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54288.11-54294.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[25]_TMR_0  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_0),
    .CK(sys_clk),
    .D(N_427_TMR_0),
    .Q(dsp_join_kb_27_TMR_0[25]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54288.11-54294.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[25]_TMR_1  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_1),
    .CK(sys_clk),
    .D(N_427_TMR_1),
    .Q(dsp_join_kb_27_TMR_1[25]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54288.11-54294.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[25]_TMR_2  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_2),
    .CK(sys_clk),
    .D(N_427_TMR_2),
    .Q(dsp_join_kb_27_TMR_2[25]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54295.11-54301.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[26]_TMR_0  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_0),
    .CK(sys_clk),
    .D(N_428_TMR_0),
    .Q(dsp_join_kb_27_TMR_0[26]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54295.11-54301.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[26]_TMR_1  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_1),
    .CK(sys_clk),
    .D(N_428_TMR_1),
    .Q(dsp_join_kb_27_TMR_1[26]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54295.11-54301.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[26]_TMR_2  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_2),
    .CK(sys_clk),
    .D(N_428_TMR_2),
    .Q(dsp_join_kb_27_TMR_2[26]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54302.11-54308.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[27]_TMR_0  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_0),
    .CK(sys_clk),
    .D(N_429_TMR_0),
    .Q(dsp_join_kb_27_TMR_0[27]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54302.11-54308.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[27]_TMR_1  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_1),
    .CK(sys_clk),
    .D(N_429_TMR_1),
    .Q(dsp_join_kb_27_TMR_1[27]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54302.11-54308.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[27]_TMR_2  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_2),
    .CK(sys_clk),
    .D(N_429_TMR_2),
    .Q(dsp_join_kb_27_TMR_2[27]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54309.11-54315.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[28]_TMR_0  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_0),
    .CK(sys_clk),
    .D(N_430_TMR_0),
    .Q(dsp_join_kb_27_TMR_0[28]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54309.11-54315.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[28]_TMR_1  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_1),
    .CK(sys_clk),
    .D(N_430_TMR_1),
    .Q(dsp_join_kb_27_TMR_1[28]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54309.11-54315.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[28]_TMR_2  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_2),
    .CK(sys_clk),
    .D(N_430_TMR_2),
    .Q(dsp_join_kb_27_TMR_2[28]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54316.11-54322.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[29]_TMR_0  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_0),
    .CK(sys_clk),
    .D(un5_main_basesoc_rx_phase_cry_29_0_S0_TMR_0),
    .Q(dsp_join_kb_27_TMR_0[29]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54316.11-54322.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[29]_TMR_1  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_1),
    .CK(sys_clk),
    .D(un5_main_basesoc_rx_phase_cry_29_0_S0_TMR_1),
    .Q(dsp_join_kb_27_TMR_1[29]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54316.11-54322.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[29]_TMR_2  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_2),
    .CK(sys_clk),
    .D(un5_main_basesoc_rx_phase_cry_29_0_S0_TMR_2),
    .Q(dsp_join_kb_27_TMR_2[29]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54127.11-54133.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[2]_TMR_0  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_0),
    .CK(sys_clk),
    .D(N_404_TMR_0),
    .Q(dsp_join_kb_27_TMR_0[2]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54127.11-54133.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[2]_TMR_1  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_1),
    .CK(sys_clk),
    .D(N_404_TMR_1),
    .Q(dsp_join_kb_27_TMR_1[2]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54127.11-54133.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[2]_TMR_2  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_2),
    .CK(sys_clk),
    .D(N_404_TMR_2),
    .Q(dsp_join_kb_27_TMR_2[2]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54323.11-54329.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[30]_TMR_0  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_0),
    .CK(sys_clk),
    .D(un5_main_basesoc_rx_phase_cry_29_0_S1_TMR_0),
    .Q(dsp_join_kb_27_TMR_0[30]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54323.11-54329.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[30]_TMR_1  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_1),
    .CK(sys_clk),
    .D(un5_main_basesoc_rx_phase_cry_29_0_S1_TMR_1),
    .Q(dsp_join_kb_27_TMR_1[30]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54323.11-54329.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[30]_TMR_2  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_2),
    .CK(sys_clk),
    .D(un5_main_basesoc_rx_phase_cry_29_0_S1_TMR_2),
    .Q(dsp_join_kb_27_TMR_2[30]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54134.11-54140.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[3]_TMR_0  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_0),
    .CK(sys_clk),
    .D(N_405_TMR_0),
    .Q(dsp_join_kb_27_TMR_0[3]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54134.11-54140.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[3]_TMR_1  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_1),
    .CK(sys_clk),
    .D(N_405_TMR_1),
    .Q(dsp_join_kb_27_TMR_1[3]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54134.11-54140.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[3]_TMR_2  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_2),
    .CK(sys_clk),
    .D(N_405_TMR_2),
    .Q(dsp_join_kb_27_TMR_2[3]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54141.11-54147.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[4]_TMR_0  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_0),
    .CK(sys_clk),
    .D(N_406_TMR_0),
    .Q(dsp_join_kb_27_TMR_0[4]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54141.11-54147.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[4]_TMR_1  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_1),
    .CK(sys_clk),
    .D(N_406_TMR_1),
    .Q(dsp_join_kb_27_TMR_1[4]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54141.11-54147.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[4]_TMR_2  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_2),
    .CK(sys_clk),
    .D(N_406_TMR_2),
    .Q(dsp_join_kb_27_TMR_2[4]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54148.11-54154.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[5]_TMR_0  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_0),
    .CK(sys_clk),
    .D(N_407_TMR_0),
    .Q(dsp_join_kb_27_TMR_0[5]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54148.11-54154.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[5]_TMR_1  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_1),
    .CK(sys_clk),
    .D(N_407_TMR_1),
    .Q(dsp_join_kb_27_TMR_1[5]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54148.11-54154.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[5]_TMR_2  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_2),
    .CK(sys_clk),
    .D(N_407_TMR_2),
    .Q(dsp_join_kb_27_TMR_2[5]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54155.11-54161.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[6]_TMR_0  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_0),
    .CK(sys_clk),
    .D(N_408_TMR_0),
    .Q(dsp_join_kb_27_TMR_0[6]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54155.11-54161.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[6]_TMR_1  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_1),
    .CK(sys_clk),
    .D(N_408_TMR_1),
    .Q(dsp_join_kb_27_TMR_1[6]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54155.11-54161.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[6]_TMR_2  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_2),
    .CK(sys_clk),
    .D(N_408_TMR_2),
    .Q(dsp_join_kb_27_TMR_2[6]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54162.11-54168.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[7]_TMR_0  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_0),
    .CK(sys_clk),
    .D(N_409_TMR_0),
    .Q(dsp_join_kb_27_TMR_0[7]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54162.11-54168.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[7]_TMR_1  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_1),
    .CK(sys_clk),
    .D(N_409_TMR_1),
    .Q(dsp_join_kb_27_TMR_1[7]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54162.11-54168.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[7]_TMR_2  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_2),
    .CK(sys_clk),
    .D(N_409_TMR_2),
    .Q(dsp_join_kb_27_TMR_2[7]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54169.11-54175.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[8]_TMR_0  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_0),
    .CK(sys_clk),
    .D(N_410_TMR_0),
    .Q(dsp_join_kb_27_TMR_0[8]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54169.11-54175.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[8]_TMR_1  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_1),
    .CK(sys_clk),
    .D(N_410_TMR_1),
    .Q(dsp_join_kb_27_TMR_1[8]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54169.11-54175.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[8]_TMR_2  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_2),
    .CK(sys_clk),
    .D(N_410_TMR_2),
    .Q(dsp_join_kb_27_TMR_2[8]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54176.11-54182.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[9]_TMR_0  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_0),
    .CK(sys_clk),
    .D(N_411_TMR_0),
    .Q(dsp_join_kb_27_TMR_0[9]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54176.11-54182.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[9]_TMR_1  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_1),
    .CK(sys_clk),
    .D(N_411_TMR_1),
    .Q(dsp_join_kb_27_TMR_1[9]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54176.11-54182.2" *)
  FD1P3IX \main_basesoc_rx_phase_mod[9]_TMR_2  (
    .CD(builder_basesoc_rs232phyrx_state_i_TMR_2),
    .CK(sys_clk),
    .D(N_411_TMR_2),
    .Q(dsp_join_kb_27_TMR_2[9]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56058.8-56064.2" *)
  LUT4 \main_basesoc_rx_phase_mod_RNO_cZ[0]_TMR_0  (
    .A(builder_basesoc_rs232phyrx_state_TMR_0),
    .B(dsp_join_kb_27_TMR_0[0]),
    .C(GND_0),
    .D(GND_0),
    .Z(main_basesoc_rx_phase_mod_RNO_TMR_0)
  );
  defparam \main_basesoc_rx_phase_mod_RNO_cZ[0]_TMR_0 .INIT = "0x2222";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56058.8-56064.2" *)
  LUT4 \main_basesoc_rx_phase_mod_RNO_cZ[0]_TMR_1  (
    .A(builder_basesoc_rs232phyrx_state_TMR_1),
    .B(dsp_join_kb_27_TMR_1[0]),
    .C(GND_0),
    .D(GND_0),
    .Z(main_basesoc_rx_phase_mod_RNO_TMR_1)
  );
  defparam \main_basesoc_rx_phase_mod_RNO_cZ[0]_TMR_1 .INIT = "0x2222";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56058.8-56064.2" *)
  LUT4 \main_basesoc_rx_phase_mod_RNO_cZ[0]_TMR_2  (
    .A(builder_basesoc_rs232phyrx_state_TMR_2),
    .B(dsp_join_kb_27_TMR_2[0]),
    .C(GND_0),
    .D(GND_0),
    .Z(main_basesoc_rx_phase_mod_RNO_TMR_2)
  );
  defparam \main_basesoc_rx_phase_mod_RNO_cZ[0]_TMR_2 .INIT = "0x2222";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54106.11-54112.2" *)
  FD1P3IX main_basesoc_rx_rx_d_reg_TMR_0 (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(builder_regs1_TMR_0),
    .Q(main_basesoc_rx_rx_d_TMR_0),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54106.11-54112.2" *)
  FD1P3IX main_basesoc_rx_rx_d_reg_TMR_1 (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(builder_regs1_TMR_1),
    .Q(main_basesoc_rx_rx_d_TMR_1),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54106.11-54112.2" *)
  FD1P3IX main_basesoc_rx_rx_d_reg_TMR_2 (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(builder_regs1_TMR_2),
    .Q(main_basesoc_rx_rx_d_TMR_2),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54099.11-54105.2" *)
  FD1P3IX main_basesoc_rx_tick_reg_TMR_0 (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(main_basesoc_rx_tick_0_TMR_0),
    .Q(main_basesoc_rx_tick_TMR_0),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54099.11-54105.2" *)
  FD1P3IX main_basesoc_rx_tick_reg_TMR_1 (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(main_basesoc_rx_tick_0_TMR_1),
    .Q(main_basesoc_rx_tick_TMR_1),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54099.11-54105.2" *)
  FD1P3IX main_basesoc_rx_tick_reg_TMR_2 (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(main_basesoc_rx_tick_0_TMR_2),
    .Q(main_basesoc_rx_tick_TMR_2),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53875.11-53881.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[0]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[0]),
    .Q(main_basesoc_scratch_storage_TMR_0[0]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53875.11-53881.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[0]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[0]),
    .Q(main_basesoc_scratch_storage_TMR_1[0]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53875.11-53881.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[0]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[0]),
    .Q(main_basesoc_scratch_storage_TMR_2[0]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53945.11-53951.2" *)
  FD1P3JX \main_basesoc_scratch_storage_reg[10]_TMR_0  (
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[10]),
    .PD(sys_rst_TMR_0),
    .Q(main_basesoc_scratch_storage_TMR_0[10]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53945.11-53951.2" *)
  FD1P3JX \main_basesoc_scratch_storage_reg[10]_TMR_1  (
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[10]),
    .PD(sys_rst_TMR_1),
    .Q(main_basesoc_scratch_storage_TMR_1[10]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53945.11-53951.2" *)
  FD1P3JX \main_basesoc_scratch_storage_reg[10]_TMR_2  (
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[10]),
    .PD(sys_rst_TMR_2),
    .Q(main_basesoc_scratch_storage_TMR_2[10]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53952.11-53958.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[11]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[11]),
    .Q(main_basesoc_scratch_storage_TMR_0[11]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53952.11-53958.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[11]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[11]),
    .Q(main_basesoc_scratch_storage_TMR_1[11]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53952.11-53958.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[11]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[11]),
    .Q(main_basesoc_scratch_storage_TMR_2[11]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53959.11-53965.2" *)
  FD1P3JX \main_basesoc_scratch_storage_reg[12]_TMR_0  (
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[12]),
    .PD(sys_rst_TMR_0),
    .Q(main_basesoc_scratch_storage_TMR_0[12]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53959.11-53965.2" *)
  FD1P3JX \main_basesoc_scratch_storage_reg[12]_TMR_1  (
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[12]),
    .PD(sys_rst_TMR_1),
    .Q(main_basesoc_scratch_storage_TMR_1[12]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53959.11-53965.2" *)
  FD1P3JX \main_basesoc_scratch_storage_reg[12]_TMR_2  (
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[12]),
    .PD(sys_rst_TMR_2),
    .Q(main_basesoc_scratch_storage_TMR_2[12]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53966.11-53972.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[13]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[13]),
    .Q(main_basesoc_scratch_storage_TMR_0[13]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53966.11-53972.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[13]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[13]),
    .Q(main_basesoc_scratch_storage_TMR_1[13]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53966.11-53972.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[13]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[13]),
    .Q(main_basesoc_scratch_storage_TMR_2[13]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53973.11-53979.2" *)
  FD1P3JX \main_basesoc_scratch_storage_reg[14]_TMR_0  (
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[14]),
    .PD(sys_rst_TMR_0),
    .Q(main_basesoc_scratch_storage_TMR_0[14]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53973.11-53979.2" *)
  FD1P3JX \main_basesoc_scratch_storage_reg[14]_TMR_1  (
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[14]),
    .PD(sys_rst_TMR_1),
    .Q(main_basesoc_scratch_storage_TMR_1[14]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53973.11-53979.2" *)
  FD1P3JX \main_basesoc_scratch_storage_reg[14]_TMR_2  (
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[14]),
    .PD(sys_rst_TMR_2),
    .Q(main_basesoc_scratch_storage_TMR_2[14]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53980.11-53986.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[15]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[15]),
    .Q(main_basesoc_scratch_storage_TMR_0[15]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53980.11-53986.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[15]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[15]),
    .Q(main_basesoc_scratch_storage_TMR_1[15]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53980.11-53986.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[15]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[15]),
    .Q(main_basesoc_scratch_storage_TMR_2[15]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53987.11-53993.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[16]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[16]),
    .Q(main_basesoc_scratch_storage_TMR_0[16]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53987.11-53993.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[16]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[16]),
    .Q(main_basesoc_scratch_storage_TMR_1[16]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53987.11-53993.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[16]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[16]),
    .Q(main_basesoc_scratch_storage_TMR_2[16]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53994.11-54000.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[17]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[17]),
    .Q(main_basesoc_scratch_storage_TMR_0[17]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53994.11-54000.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[17]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[17]),
    .Q(main_basesoc_scratch_storage_TMR_1[17]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53994.11-54000.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[17]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[17]),
    .Q(main_basesoc_scratch_storage_TMR_2[17]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54001.11-54007.2" *)
  FD1P3JX \main_basesoc_scratch_storage_reg[18]_TMR_0  (
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[18]),
    .PD(sys_rst_TMR_0),
    .Q(main_basesoc_scratch_storage_TMR_0[18]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54001.11-54007.2" *)
  FD1P3JX \main_basesoc_scratch_storage_reg[18]_TMR_1  (
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[18]),
    .PD(sys_rst_TMR_1),
    .Q(main_basesoc_scratch_storage_TMR_1[18]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54001.11-54007.2" *)
  FD1P3JX \main_basesoc_scratch_storage_reg[18]_TMR_2  (
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[18]),
    .PD(sys_rst_TMR_2),
    .Q(main_basesoc_scratch_storage_TMR_2[18]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54008.11-54014.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[19]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[19]),
    .Q(main_basesoc_scratch_storage_TMR_0[19]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54008.11-54014.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[19]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[19]),
    .Q(main_basesoc_scratch_storage_TMR_1[19]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54008.11-54014.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[19]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[19]),
    .Q(main_basesoc_scratch_storage_TMR_2[19]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53882.11-53888.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[1]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[1]),
    .Q(main_basesoc_scratch_storage_TMR_0[1]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53882.11-53888.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[1]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[1]),
    .Q(main_basesoc_scratch_storage_TMR_1[1]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53882.11-53888.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[1]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[1]),
    .Q(main_basesoc_scratch_storage_TMR_2[1]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54015.11-54021.2" *)
  FD1P3JX \main_basesoc_scratch_storage_reg[20]_TMR_0  (
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[20]),
    .PD(sys_rst_TMR_0),
    .Q(main_basesoc_scratch_storage_TMR_0[20]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54015.11-54021.2" *)
  FD1P3JX \main_basesoc_scratch_storage_reg[20]_TMR_1  (
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[20]),
    .PD(sys_rst_TMR_1),
    .Q(main_basesoc_scratch_storage_TMR_1[20]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54015.11-54021.2" *)
  FD1P3JX \main_basesoc_scratch_storage_reg[20]_TMR_2  (
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[20]),
    .PD(sys_rst_TMR_2),
    .Q(main_basesoc_scratch_storage_TMR_2[20]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54022.11-54028.2" *)
  FD1P3JX \main_basesoc_scratch_storage_reg[21]_TMR_0  (
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[21]),
    .PD(sys_rst_TMR_0),
    .Q(main_basesoc_scratch_storage_TMR_0[21]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54022.11-54028.2" *)
  FD1P3JX \main_basesoc_scratch_storage_reg[21]_TMR_1  (
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[21]),
    .PD(sys_rst_TMR_1),
    .Q(main_basesoc_scratch_storage_TMR_1[21]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54022.11-54028.2" *)
  FD1P3JX \main_basesoc_scratch_storage_reg[21]_TMR_2  (
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[21]),
    .PD(sys_rst_TMR_2),
    .Q(main_basesoc_scratch_storage_TMR_2[21]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54029.11-54035.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[22]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[22]),
    .Q(main_basesoc_scratch_storage_TMR_0[22]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54029.11-54035.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[22]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[22]),
    .Q(main_basesoc_scratch_storage_TMR_1[22]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54029.11-54035.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[22]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[22]),
    .Q(main_basesoc_scratch_storage_TMR_2[22]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54036.11-54042.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[23]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[23]),
    .Q(main_basesoc_scratch_storage_TMR_0[23]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54036.11-54042.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[23]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[23]),
    .Q(main_basesoc_scratch_storage_TMR_1[23]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54036.11-54042.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[23]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[23]),
    .Q(main_basesoc_scratch_storage_TMR_2[23]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54043.11-54049.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[24]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[24]),
    .Q(main_basesoc_scratch_storage_TMR_0[24]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54043.11-54049.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[24]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[24]),
    .Q(main_basesoc_scratch_storage_TMR_1[24]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54043.11-54049.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[24]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[24]),
    .Q(main_basesoc_scratch_storage_TMR_2[24]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54050.11-54056.2" *)
  FD1P3JX \main_basesoc_scratch_storage_reg[25]_TMR_0  (
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[25]),
    .PD(sys_rst_TMR_0),
    .Q(main_basesoc_scratch_storage_TMR_0[25]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54050.11-54056.2" *)
  FD1P3JX \main_basesoc_scratch_storage_reg[25]_TMR_1  (
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[25]),
    .PD(sys_rst_TMR_1),
    .Q(main_basesoc_scratch_storage_TMR_1[25]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54050.11-54056.2" *)
  FD1P3JX \main_basesoc_scratch_storage_reg[25]_TMR_2  (
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[25]),
    .PD(sys_rst_TMR_2),
    .Q(main_basesoc_scratch_storage_TMR_2[25]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54057.11-54063.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[26]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_split_kb_0_TMR_0),
    .Q(main_basesoc_scratch_storage_TMR_0[26]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54057.11-54063.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[26]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_split_kb_0_TMR_1),
    .Q(main_basesoc_scratch_storage_TMR_1[26]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54057.11-54063.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[26]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_split_kb_0_TMR_2),
    .Q(main_basesoc_scratch_storage_TMR_2[26]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54064.11-54070.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[27]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[26]),
    .Q(main_basesoc_scratch_storage_TMR_0[27]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54064.11-54070.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[27]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[26]),
    .Q(main_basesoc_scratch_storage_TMR_1[27]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54064.11-54070.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[27]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[26]),
    .Q(main_basesoc_scratch_storage_TMR_2[27]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54071.11-54077.2" *)
  FD1P3JX \main_basesoc_scratch_storage_reg[28]_TMR_0  (
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[27]),
    .PD(sys_rst_TMR_0),
    .Q(main_basesoc_scratch_storage_TMR_0[28]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54071.11-54077.2" *)
  FD1P3JX \main_basesoc_scratch_storage_reg[28]_TMR_1  (
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[27]),
    .PD(sys_rst_TMR_1),
    .Q(main_basesoc_scratch_storage_TMR_1[28]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54071.11-54077.2" *)
  FD1P3JX \main_basesoc_scratch_storage_reg[28]_TMR_2  (
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[27]),
    .PD(sys_rst_TMR_2),
    .Q(main_basesoc_scratch_storage_TMR_2[28]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54078.11-54084.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[29]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[28]),
    .Q(main_basesoc_scratch_storage_TMR_0[29]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54078.11-54084.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[29]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[28]),
    .Q(main_basesoc_scratch_storage_TMR_1[29]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54078.11-54084.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[29]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[28]),
    .Q(main_basesoc_scratch_storage_TMR_2[29]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53889.11-53895.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[2]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[2]),
    .Q(main_basesoc_scratch_storage_TMR_0[2]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53889.11-53895.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[2]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[2]),
    .Q(main_basesoc_scratch_storage_TMR_1[2]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53889.11-53895.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[2]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[2]),
    .Q(main_basesoc_scratch_storage_TMR_2[2]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54085.11-54091.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[30]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[29]),
    .Q(main_basesoc_scratch_storage_TMR_0[30]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54085.11-54091.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[30]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[29]),
    .Q(main_basesoc_scratch_storage_TMR_1[30]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54085.11-54091.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[30]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[29]),
    .Q(main_basesoc_scratch_storage_TMR_2[30]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54092.11-54098.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[31]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[30]),
    .Q(main_basesoc_scratch_storage_TMR_0[31]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54092.11-54098.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[31]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[30]),
    .Q(main_basesoc_scratch_storage_TMR_1[31]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:54092.11-54098.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[31]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[30]),
    .Q(main_basesoc_scratch_storage_TMR_2[31]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53896.11-53902.2" *)
  FD1P3JX \main_basesoc_scratch_storage_reg[3]_TMR_0  (
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[3]),
    .PD(sys_rst_TMR_0),
    .Q(main_basesoc_scratch_storage_TMR_0[3]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53896.11-53902.2" *)
  FD1P3JX \main_basesoc_scratch_storage_reg[3]_TMR_1  (
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[3]),
    .PD(sys_rst_TMR_1),
    .Q(main_basesoc_scratch_storage_TMR_1[3]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53896.11-53902.2" *)
  FD1P3JX \main_basesoc_scratch_storage_reg[3]_TMR_2  (
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[3]),
    .PD(sys_rst_TMR_2),
    .Q(main_basesoc_scratch_storage_TMR_2[3]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53903.11-53909.2" *)
  FD1P3JX \main_basesoc_scratch_storage_reg[4]_TMR_0  (
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[4]),
    .PD(sys_rst_TMR_0),
    .Q(main_basesoc_scratch_storage_TMR_0[4]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53903.11-53909.2" *)
  FD1P3JX \main_basesoc_scratch_storage_reg[4]_TMR_1  (
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[4]),
    .PD(sys_rst_TMR_1),
    .Q(main_basesoc_scratch_storage_TMR_1[4]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53903.11-53909.2" *)
  FD1P3JX \main_basesoc_scratch_storage_reg[4]_TMR_2  (
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[4]),
    .PD(sys_rst_TMR_2),
    .Q(main_basesoc_scratch_storage_TMR_2[4]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53910.11-53916.2" *)
  FD1P3JX \main_basesoc_scratch_storage_reg[5]_TMR_0  (
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[5]),
    .PD(sys_rst_TMR_0),
    .Q(main_basesoc_scratch_storage_TMR_0[5]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53910.11-53916.2" *)
  FD1P3JX \main_basesoc_scratch_storage_reg[5]_TMR_1  (
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[5]),
    .PD(sys_rst_TMR_1),
    .Q(main_basesoc_scratch_storage_TMR_1[5]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53910.11-53916.2" *)
  FD1P3JX \main_basesoc_scratch_storage_reg[5]_TMR_2  (
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[5]),
    .PD(sys_rst_TMR_2),
    .Q(main_basesoc_scratch_storage_TMR_2[5]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53917.11-53923.2" *)
  FD1P3JX \main_basesoc_scratch_storage_reg[6]_TMR_0  (
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[6]),
    .PD(sys_rst_TMR_0),
    .Q(main_basesoc_scratch_storage_TMR_0[6]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53917.11-53923.2" *)
  FD1P3JX \main_basesoc_scratch_storage_reg[6]_TMR_1  (
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[6]),
    .PD(sys_rst_TMR_1),
    .Q(main_basesoc_scratch_storage_TMR_1[6]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53917.11-53923.2" *)
  FD1P3JX \main_basesoc_scratch_storage_reg[6]_TMR_2  (
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[6]),
    .PD(sys_rst_TMR_2),
    .Q(main_basesoc_scratch_storage_TMR_2[6]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53924.11-53930.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[7]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[7]),
    .Q(main_basesoc_scratch_storage_TMR_0[7]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53924.11-53930.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[7]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[7]),
    .Q(main_basesoc_scratch_storage_TMR_1[7]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53924.11-53930.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[7]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[7]),
    .Q(main_basesoc_scratch_storage_TMR_2[7]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53931.11-53937.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[8]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[8]),
    .Q(main_basesoc_scratch_storage_TMR_0[8]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53931.11-53937.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[8]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[8]),
    .Q(main_basesoc_scratch_storage_TMR_1[8]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53931.11-53937.2" *)
  FD1P3IX \main_basesoc_scratch_storage_reg[8]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[8]),
    .Q(main_basesoc_scratch_storage_TMR_2[8]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53938.11-53944.2" *)
  FD1P3JX \main_basesoc_scratch_storage_reg[9]_TMR_0  (
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[9]),
    .PD(sys_rst_TMR_0),
    .Q(main_basesoc_scratch_storage_TMR_0[9]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53938.11-53944.2" *)
  FD1P3JX \main_basesoc_scratch_storage_reg[9]_TMR_1  (
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[9]),
    .PD(sys_rst_TMR_1),
    .Q(main_basesoc_scratch_storage_TMR_1[9]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53938.11-53944.2" *)
  FD1P3JX \main_basesoc_scratch_storage_reg[9]_TMR_2  (
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[9]),
    .PD(sys_rst_TMR_2),
    .Q(main_basesoc_scratch_storage_TMR_2[9]),
    .SP(builder_csr_bankarray_csrbank0_scratch0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53868.11-53874.2" *)
  FD1P3IX main_basesoc_timer_en_storage_reg_TMR_0 (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[0]),
    .Q(main_basesoc_timer_en_storage_TMR_0),
    .SP(builder_csr_bankarray_csrbank2_en0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53868.11-53874.2" *)
  FD1P3IX main_basesoc_timer_en_storage_reg_TMR_1 (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[0]),
    .Q(main_basesoc_timer_en_storage_TMR_1),
    .SP(builder_csr_bankarray_csrbank2_en0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53868.11-53874.2" *)
  FD1P3IX main_basesoc_timer_en_storage_reg_TMR_2 (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[0]),
    .Q(main_basesoc_timer_en_storage_TMR_2),
    .SP(builder_csr_bankarray_csrbank2_en0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53861.11-53867.2" *)
  FD1P3IX main_basesoc_timer_enable_storage_reg_TMR_0 (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[0]),
    .Q(main_basesoc_timer_enable_storage_TMR_0),
    .SP(builder_csr_bankarray_csrbank2_ev_enable0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53861.11-53867.2" *)
  FD1P3IX main_basesoc_timer_enable_storage_reg_TMR_1 (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[0]),
    .Q(main_basesoc_timer_enable_storage_TMR_1),
    .SP(builder_csr_bankarray_csrbank2_ev_enable0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53861.11-53867.2" *)
  FD1P3IX main_basesoc_timer_enable_storage_reg_TMR_2 (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[0]),
    .Q(main_basesoc_timer_enable_storage_TMR_2),
    .SP(builder_csr_bankarray_csrbank2_ev_enable0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53749.11-53755.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_0_mod[0]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_timer_load_storage_0_mod_RNO_TMR_0),
    .Q(dsp_join_kb_TMR_0[0]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53749.11-53755.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_0_mod[0]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_timer_load_storage_0_mod_RNO_TMR_1),
    .Q(dsp_join_kb_TMR_1[0]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53749.11-53755.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_0_mod[0]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_timer_load_storage_0_mod_RNO_TMR_2),
    .Q(dsp_join_kb_TMR_2[0]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53784.11-53790.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_0_mod[10]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[10]),
    .Q(dsp_join_kb_TMR_0[10]),
    .SP(N_443_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53784.11-53790.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_0_mod[10]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[10]),
    .Q(dsp_join_kb_TMR_1[10]),
    .SP(N_443_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53784.11-53790.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_0_mod[10]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[10]),
    .Q(dsp_join_kb_TMR_2[10]),
    .SP(N_443_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53791.11-53797.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_0_mod[12]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[12]),
    .Q(dsp_join_kb_TMR_0[12]),
    .SP(N_443_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53791.11-53797.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_0_mod[12]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[12]),
    .Q(dsp_join_kb_TMR_1[12]),
    .SP(N_443_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53791.11-53797.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_0_mod[12]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[12]),
    .Q(dsp_join_kb_TMR_2[12]),
    .SP(N_443_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53798.11-53804.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_0_mod[14]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[14]),
    .Q(dsp_join_kb_TMR_0[14]),
    .SP(N_443_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53798.11-53804.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_0_mod[14]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[14]),
    .Q(dsp_join_kb_TMR_1[14]),
    .SP(N_443_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53798.11-53804.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_0_mod[14]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[14]),
    .Q(dsp_join_kb_TMR_2[14]),
    .SP(N_443_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53805.11-53811.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_0_mod[16]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[16]),
    .Q(dsp_join_kb_TMR_0[16]),
    .SP(N_443_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53805.11-53811.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_0_mod[16]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[16]),
    .Q(dsp_join_kb_TMR_1[16]),
    .SP(N_443_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53805.11-53811.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_0_mod[16]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[16]),
    .Q(dsp_join_kb_TMR_2[16]),
    .SP(N_443_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53812.11-53818.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_0_mod[18]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[18]),
    .Q(dsp_join_kb_TMR_0[18]),
    .SP(N_443_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53812.11-53818.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_0_mod[18]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[18]),
    .Q(dsp_join_kb_TMR_1[18]),
    .SP(N_443_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53812.11-53818.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_0_mod[18]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[18]),
    .Q(dsp_join_kb_TMR_2[18]),
    .SP(N_443_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53819.11-53825.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_0_mod[20]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[20]),
    .Q(dsp_join_kb_TMR_0[20]),
    .SP(N_443_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53819.11-53825.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_0_mod[20]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[20]),
    .Q(dsp_join_kb_TMR_1[20]),
    .SP(N_443_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53819.11-53825.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_0_mod[20]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[20]),
    .Q(dsp_join_kb_TMR_2[20]),
    .SP(N_443_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53826.11-53832.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_0_mod[22]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[22]),
    .Q(dsp_join_kb_TMR_0[22]),
    .SP(N_443_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53826.11-53832.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_0_mod[22]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[22]),
    .Q(dsp_join_kb_TMR_1[22]),
    .SP(N_443_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53826.11-53832.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_0_mod[22]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[22]),
    .Q(dsp_join_kb_TMR_2[22]),
    .SP(N_443_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53833.11-53839.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_0_mod[24]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[24]),
    .Q(dsp_join_kb_TMR_0[24]),
    .SP(N_443_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53833.11-53839.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_0_mod[24]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[24]),
    .Q(dsp_join_kb_TMR_1[24]),
    .SP(N_443_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53833.11-53839.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_0_mod[24]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[24]),
    .Q(dsp_join_kb_TMR_2[24]),
    .SP(N_443_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53840.11-53846.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_0_mod[26]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_split_kb_0_TMR_0),
    .Q(dsp_split_kb_1_TMR_0),
    .SP(N_443_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53840.11-53846.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_0_mod[26]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_split_kb_0_TMR_1),
    .Q(dsp_split_kb_1_TMR_1),
    .SP(N_443_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53840.11-53846.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_0_mod[26]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_split_kb_0_TMR_2),
    .Q(dsp_split_kb_1_TMR_2),
    .SP(N_443_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53847.11-53853.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_0_mod[28]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[27]),
    .Q(dsp_join_kb_TMR_0[27]),
    .SP(N_443_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53847.11-53853.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_0_mod[28]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[27]),
    .Q(dsp_join_kb_TMR_1[27]),
    .SP(N_443_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53847.11-53853.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_0_mod[28]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[27]),
    .Q(dsp_join_kb_TMR_2[27]),
    .SP(N_443_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53756.11-53762.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_0_mod[2]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[2]),
    .Q(dsp_join_kb_TMR_0[2]),
    .SP(N_443_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53756.11-53762.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_0_mod[2]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[2]),
    .Q(dsp_join_kb_TMR_1[2]),
    .SP(N_443_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53756.11-53762.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_0_mod[2]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[2]),
    .Q(dsp_join_kb_TMR_2[2]),
    .SP(N_443_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53854.11-53860.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_0_mod[30]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[29]),
    .Q(dsp_join_kb_TMR_0[29]),
    .SP(N_443_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53854.11-53860.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_0_mod[30]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[29]),
    .Q(dsp_join_kb_TMR_1[29]),
    .SP(N_443_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53854.11-53860.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_0_mod[30]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[29]),
    .Q(dsp_join_kb_TMR_2[29]),
    .SP(N_443_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53763.11-53769.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_0_mod[4]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[4]),
    .Q(dsp_join_kb_TMR_0[4]),
    .SP(N_443_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53763.11-53769.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_0_mod[4]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[4]),
    .Q(dsp_join_kb_TMR_1[4]),
    .SP(N_443_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53763.11-53769.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_0_mod[4]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[4]),
    .Q(dsp_join_kb_TMR_2[4]),
    .SP(N_443_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53770.11-53776.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_0_mod[6]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[6]),
    .Q(dsp_join_kb_TMR_0[6]),
    .SP(N_443_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53770.11-53776.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_0_mod[6]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[6]),
    .Q(dsp_join_kb_TMR_1[6]),
    .SP(N_443_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53770.11-53776.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_0_mod[6]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[6]),
    .Q(dsp_join_kb_TMR_2[6]),
    .SP(N_443_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53777.11-53783.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_0_mod[8]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[8]),
    .Q(dsp_join_kb_TMR_0[8]),
    .SP(N_443_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53777.11-53783.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_0_mod[8]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[8]),
    .Q(dsp_join_kb_TMR_1[8]),
    .SP(N_443_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53777.11-53783.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_0_mod[8]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[8]),
    .Q(dsp_join_kb_TMR_2[8]),
    .SP(N_443_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55870.8-55876.2" *)
  LUT4 \main_basesoc_timer_load_storage_0_mod_RNO_cZ[0]_TMR_0  (
    .A(N_443_TMR_0),
    .B(sys_rst_TMR_0),
    .C(dsp_join_kb_TMR_0[0]),
    .D(dsp_join_kb_0_TMR_0[0]),
    .Z(main_basesoc_timer_load_storage_0_mod_RNO_TMR_0)
  );
  defparam \main_basesoc_timer_load_storage_0_mod_RNO_cZ[0]_TMR_0 .INIT = "0x3210";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55870.8-55876.2" *)
  LUT4 \main_basesoc_timer_load_storage_0_mod_RNO_cZ[0]_TMR_1  (
    .A(N_443_TMR_1),
    .B(sys_rst_TMR_1),
    .C(dsp_join_kb_TMR_1[0]),
    .D(dsp_join_kb_0_TMR_1[0]),
    .Z(main_basesoc_timer_load_storage_0_mod_RNO_TMR_1)
  );
  defparam \main_basesoc_timer_load_storage_0_mod_RNO_cZ[0]_TMR_1 .INIT = "0x3210";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55870.8-55876.2" *)
  LUT4 \main_basesoc_timer_load_storage_0_mod_RNO_cZ[0]_TMR_2  (
    .A(N_443_TMR_2),
    .B(sys_rst_TMR_2),
    .C(dsp_join_kb_TMR_2[0]),
    .D(dsp_join_kb_0_TMR_2[0]),
    .Z(main_basesoc_timer_load_storage_0_mod_RNO_TMR_2)
  );
  defparam \main_basesoc_timer_load_storage_0_mod_RNO_cZ[0]_TMR_2 .INIT = "0x3210";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53672.11-53678.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_mod[11]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[11]),
    .Q(dsp_join_kb_TMR_0[11]),
    .SP(N_443_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53672.11-53678.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_mod[11]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[11]),
    .Q(dsp_join_kb_TMR_1[11]),
    .SP(N_443_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53672.11-53678.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_mod[11]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[11]),
    .Q(dsp_join_kb_TMR_2[11]),
    .SP(N_443_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53679.11-53685.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_mod[13]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[13]),
    .Q(dsp_join_kb_TMR_0[13]),
    .SP(N_443_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53679.11-53685.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_mod[13]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[13]),
    .Q(dsp_join_kb_TMR_1[13]),
    .SP(N_443_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53679.11-53685.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_mod[13]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[13]),
    .Q(dsp_join_kb_TMR_2[13]),
    .SP(N_443_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53686.11-53692.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_mod[15]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[15]),
    .Q(dsp_join_kb_TMR_0[15]),
    .SP(N_443_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53686.11-53692.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_mod[15]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[15]),
    .Q(dsp_join_kb_TMR_1[15]),
    .SP(N_443_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53686.11-53692.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_mod[15]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[15]),
    .Q(dsp_join_kb_TMR_2[15]),
    .SP(N_443_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53693.11-53699.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_mod[17]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[17]),
    .Q(dsp_join_kb_TMR_0[17]),
    .SP(N_443_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53693.11-53699.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_mod[17]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[17]),
    .Q(dsp_join_kb_TMR_1[17]),
    .SP(N_443_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53693.11-53699.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_mod[17]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[17]),
    .Q(dsp_join_kb_TMR_2[17]),
    .SP(N_443_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53700.11-53706.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_mod[19]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[19]),
    .Q(dsp_join_kb_TMR_0[19]),
    .SP(N_443_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53700.11-53706.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_mod[19]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[19]),
    .Q(dsp_join_kb_TMR_1[19]),
    .SP(N_443_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53700.11-53706.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_mod[19]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[19]),
    .Q(dsp_join_kb_TMR_2[19]),
    .SP(N_443_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53637.11-53643.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_mod[1]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[1]),
    .Q(dsp_join_kb_TMR_0[1]),
    .SP(N_443_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53637.11-53643.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_mod[1]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[1]),
    .Q(dsp_join_kb_TMR_1[1]),
    .SP(N_443_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53637.11-53643.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_mod[1]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[1]),
    .Q(dsp_join_kb_TMR_2[1]),
    .SP(N_443_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53707.11-53713.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_mod[21]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[21]),
    .Q(dsp_join_kb_TMR_0[21]),
    .SP(N_443_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53707.11-53713.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_mod[21]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[21]),
    .Q(dsp_join_kb_TMR_1[21]),
    .SP(N_443_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53707.11-53713.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_mod[21]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[21]),
    .Q(dsp_join_kb_TMR_2[21]),
    .SP(N_443_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53714.11-53720.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_mod[23]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[23]),
    .Q(dsp_join_kb_TMR_0[23]),
    .SP(N_443_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53714.11-53720.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_mod[23]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[23]),
    .Q(dsp_join_kb_TMR_1[23]),
    .SP(N_443_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53714.11-53720.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_mod[23]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[23]),
    .Q(dsp_join_kb_TMR_2[23]),
    .SP(N_443_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53721.11-53727.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_mod[25]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[25]),
    .Q(dsp_join_kb_TMR_0[25]),
    .SP(N_443_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53721.11-53727.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_mod[25]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[25]),
    .Q(dsp_join_kb_TMR_1[25]),
    .SP(N_443_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53721.11-53727.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_mod[25]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[25]),
    .Q(dsp_join_kb_TMR_2[25]),
    .SP(N_443_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53728.11-53734.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_mod[27]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[26]),
    .Q(dsp_join_kb_TMR_0[26]),
    .SP(N_443_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53728.11-53734.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_mod[27]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[26]),
    .Q(dsp_join_kb_TMR_1[26]),
    .SP(N_443_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53728.11-53734.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_mod[27]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[26]),
    .Q(dsp_join_kb_TMR_2[26]),
    .SP(N_443_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53735.11-53741.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_mod[29]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[28]),
    .Q(dsp_join_kb_TMR_0[28]),
    .SP(N_443_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53735.11-53741.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_mod[29]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[28]),
    .Q(dsp_join_kb_TMR_1[28]),
    .SP(N_443_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53735.11-53741.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_mod[29]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[28]),
    .Q(dsp_join_kb_TMR_2[28]),
    .SP(N_443_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53742.11-53748.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_mod[31]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[30]),
    .Q(dsp_join_kb_TMR_0[30]),
    .SP(N_443_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53742.11-53748.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_mod[31]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[30]),
    .Q(dsp_join_kb_TMR_1[30]),
    .SP(N_443_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53742.11-53748.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_mod[31]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[30]),
    .Q(dsp_join_kb_TMR_2[30]),
    .SP(N_443_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53644.11-53650.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_mod[3]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[3]),
    .Q(dsp_join_kb_TMR_0[3]),
    .SP(N_443_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53644.11-53650.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_mod[3]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[3]),
    .Q(dsp_join_kb_TMR_1[3]),
    .SP(N_443_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53644.11-53650.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_mod[3]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[3]),
    .Q(dsp_join_kb_TMR_2[3]),
    .SP(N_443_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53651.11-53657.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_mod[5]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[5]),
    .Q(dsp_join_kb_TMR_0[5]),
    .SP(N_443_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53651.11-53657.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_mod[5]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[5]),
    .Q(dsp_join_kb_TMR_1[5]),
    .SP(N_443_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53651.11-53657.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_mod[5]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[5]),
    .Q(dsp_join_kb_TMR_2[5]),
    .SP(N_443_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53658.11-53664.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_mod[7]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[7]),
    .Q(dsp_join_kb_TMR_0[7]),
    .SP(N_443_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53658.11-53664.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_mod[7]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[7]),
    .Q(dsp_join_kb_TMR_1[7]),
    .SP(N_443_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53658.11-53664.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_mod[7]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[7]),
    .Q(dsp_join_kb_TMR_2[7]),
    .SP(N_443_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53665.11-53671.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_mod[9]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[9]),
    .Q(dsp_join_kb_TMR_0[9]),
    .SP(N_443_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53665.11-53671.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_mod[9]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[9]),
    .Q(dsp_join_kb_TMR_1[9]),
    .SP(N_443_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53665.11-53671.2" *)
  FD1P3IX \main_basesoc_timer_load_storage_mod[9]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[9]),
    .Q(dsp_join_kb_TMR_2[9]),
    .SP(N_443_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53630.11-53636.2" *)
  FD1P3IX main_basesoc_timer_pending_r_reg_TMR_0 (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[0]),
    .Q(main_basesoc_timer_pending_r_TMR_0),
    .SP(builder_csr_bankarray_csrbank2_ev_pending_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53630.11-53636.2" *)
  FD1P3IX main_basesoc_timer_pending_r_reg_TMR_1 (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[0]),
    .Q(main_basesoc_timer_pending_r_TMR_1),
    .SP(builder_csr_bankarray_csrbank2_ev_pending_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53630.11-53636.2" *)
  FD1P3IX main_basesoc_timer_pending_r_reg_TMR_2 (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[0]),
    .Q(main_basesoc_timer_pending_r_TMR_2),
    .SP(builder_csr_bankarray_csrbank2_ev_pending_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53623.11-53629.2" *)
  FD1P3IX main_basesoc_timer_pending_re_reg_TMR_0 (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_timer_pending_r_0_sqmuxa_TMR_0),
    .Q(main_basesoc_timer_pending_re_TMR_0),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53623.11-53629.2" *)
  FD1P3IX main_basesoc_timer_pending_re_reg_TMR_1 (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_timer_pending_r_0_sqmuxa_TMR_1),
    .Q(main_basesoc_timer_pending_re_TMR_1),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53623.11-53629.2" *)
  FD1P3IX main_basesoc_timer_pending_re_reg_TMR_2 (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_timer_pending_r_0_sqmuxa_TMR_2),
    .Q(main_basesoc_timer_pending_re_TMR_2),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53399.11-53405.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[0]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[0]),
    .Q(main_basesoc_timer_reload_storage_TMR_0[0]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53399.11-53405.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[0]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[0]),
    .Q(main_basesoc_timer_reload_storage_TMR_1[0]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53399.11-53405.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[0]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[0]),
    .Q(main_basesoc_timer_reload_storage_TMR_2[0]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53469.11-53475.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[10]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[10]),
    .Q(main_basesoc_timer_reload_storage_TMR_0[10]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53469.11-53475.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[10]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[10]),
    .Q(main_basesoc_timer_reload_storage_TMR_1[10]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53469.11-53475.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[10]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[10]),
    .Q(main_basesoc_timer_reload_storage_TMR_2[10]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53476.11-53482.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[11]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[11]),
    .Q(main_basesoc_timer_reload_storage_TMR_0[11]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53476.11-53482.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[11]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[11]),
    .Q(main_basesoc_timer_reload_storage_TMR_1[11]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53476.11-53482.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[11]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[11]),
    .Q(main_basesoc_timer_reload_storage_TMR_2[11]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53483.11-53489.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[12]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[12]),
    .Q(main_basesoc_timer_reload_storage_TMR_0[12]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53483.11-53489.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[12]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[12]),
    .Q(main_basesoc_timer_reload_storage_TMR_1[12]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53483.11-53489.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[12]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[12]),
    .Q(main_basesoc_timer_reload_storage_TMR_2[12]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53490.11-53496.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[13]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[13]),
    .Q(main_basesoc_timer_reload_storage_TMR_0[13]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53490.11-53496.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[13]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[13]),
    .Q(main_basesoc_timer_reload_storage_TMR_1[13]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53490.11-53496.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[13]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[13]),
    .Q(main_basesoc_timer_reload_storage_TMR_2[13]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53497.11-53503.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[14]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[14]),
    .Q(main_basesoc_timer_reload_storage_TMR_0[14]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53497.11-53503.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[14]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[14]),
    .Q(main_basesoc_timer_reload_storage_TMR_1[14]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53497.11-53503.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[14]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[14]),
    .Q(main_basesoc_timer_reload_storage_TMR_2[14]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53504.11-53510.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[15]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[15]),
    .Q(main_basesoc_timer_reload_storage_TMR_0[15]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53504.11-53510.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[15]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[15]),
    .Q(main_basesoc_timer_reload_storage_TMR_1[15]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53504.11-53510.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[15]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[15]),
    .Q(main_basesoc_timer_reload_storage_TMR_2[15]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53511.11-53517.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[16]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[16]),
    .Q(main_basesoc_timer_reload_storage_TMR_0[16]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53511.11-53517.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[16]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[16]),
    .Q(main_basesoc_timer_reload_storage_TMR_1[16]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53511.11-53517.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[16]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[16]),
    .Q(main_basesoc_timer_reload_storage_TMR_2[16]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53518.11-53524.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[17]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[17]),
    .Q(main_basesoc_timer_reload_storage_TMR_0[17]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53518.11-53524.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[17]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[17]),
    .Q(main_basesoc_timer_reload_storage_TMR_1[17]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53518.11-53524.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[17]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[17]),
    .Q(main_basesoc_timer_reload_storage_TMR_2[17]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53525.11-53531.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[18]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[18]),
    .Q(main_basesoc_timer_reload_storage_TMR_0[18]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53525.11-53531.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[18]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[18]),
    .Q(main_basesoc_timer_reload_storage_TMR_1[18]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53525.11-53531.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[18]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[18]),
    .Q(main_basesoc_timer_reload_storage_TMR_2[18]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53532.11-53538.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[19]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[19]),
    .Q(main_basesoc_timer_reload_storage_TMR_0[19]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53532.11-53538.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[19]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[19]),
    .Q(main_basesoc_timer_reload_storage_TMR_1[19]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53532.11-53538.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[19]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[19]),
    .Q(main_basesoc_timer_reload_storage_TMR_2[19]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53406.11-53412.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[1]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[1]),
    .Q(main_basesoc_timer_reload_storage_TMR_0[1]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53406.11-53412.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[1]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[1]),
    .Q(main_basesoc_timer_reload_storage_TMR_1[1]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53406.11-53412.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[1]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[1]),
    .Q(main_basesoc_timer_reload_storage_TMR_2[1]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53539.11-53545.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[20]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[20]),
    .Q(main_basesoc_timer_reload_storage_TMR_0[20]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53539.11-53545.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[20]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[20]),
    .Q(main_basesoc_timer_reload_storage_TMR_1[20]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53539.11-53545.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[20]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[20]),
    .Q(main_basesoc_timer_reload_storage_TMR_2[20]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53546.11-53552.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[21]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[21]),
    .Q(main_basesoc_timer_reload_storage_TMR_0[21]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53546.11-53552.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[21]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[21]),
    .Q(main_basesoc_timer_reload_storage_TMR_1[21]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53546.11-53552.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[21]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[21]),
    .Q(main_basesoc_timer_reload_storage_TMR_2[21]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53553.11-53559.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[22]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[22]),
    .Q(main_basesoc_timer_reload_storage_TMR_0[22]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53553.11-53559.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[22]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[22]),
    .Q(main_basesoc_timer_reload_storage_TMR_1[22]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53553.11-53559.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[22]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[22]),
    .Q(main_basesoc_timer_reload_storage_TMR_2[22]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53560.11-53566.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[23]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[23]),
    .Q(main_basesoc_timer_reload_storage_TMR_0[23]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53560.11-53566.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[23]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[23]),
    .Q(main_basesoc_timer_reload_storage_TMR_1[23]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53560.11-53566.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[23]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[23]),
    .Q(main_basesoc_timer_reload_storage_TMR_2[23]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53567.11-53573.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[24]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[24]),
    .Q(main_basesoc_timer_reload_storage_TMR_0[24]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53567.11-53573.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[24]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[24]),
    .Q(main_basesoc_timer_reload_storage_TMR_1[24]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53567.11-53573.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[24]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[24]),
    .Q(main_basesoc_timer_reload_storage_TMR_2[24]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53574.11-53580.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[25]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[25]),
    .Q(main_basesoc_timer_reload_storage_TMR_0[25]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53574.11-53580.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[25]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[25]),
    .Q(main_basesoc_timer_reload_storage_TMR_1[25]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53574.11-53580.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[25]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[25]),
    .Q(main_basesoc_timer_reload_storage_TMR_2[25]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53581.11-53587.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[26]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_split_kb_0_TMR_0),
    .Q(main_basesoc_timer_reload_storage_TMR_0[26]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53581.11-53587.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[26]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_split_kb_0_TMR_1),
    .Q(main_basesoc_timer_reload_storage_TMR_1[26]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53581.11-53587.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[26]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_split_kb_0_TMR_2),
    .Q(main_basesoc_timer_reload_storage_TMR_2[26]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53588.11-53594.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[27]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[26]),
    .Q(main_basesoc_timer_reload_storage_TMR_0[27]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53588.11-53594.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[27]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[26]),
    .Q(main_basesoc_timer_reload_storage_TMR_1[27]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53588.11-53594.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[27]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[26]),
    .Q(main_basesoc_timer_reload_storage_TMR_2[27]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53595.11-53601.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[28]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[27]),
    .Q(main_basesoc_timer_reload_storage_TMR_0[28]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53595.11-53601.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[28]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[27]),
    .Q(main_basesoc_timer_reload_storage_TMR_1[28]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53595.11-53601.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[28]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[27]),
    .Q(main_basesoc_timer_reload_storage_TMR_2[28]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53602.11-53608.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[29]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[28]),
    .Q(main_basesoc_timer_reload_storage_TMR_0[29]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53602.11-53608.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[29]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[28]),
    .Q(main_basesoc_timer_reload_storage_TMR_1[29]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53602.11-53608.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[29]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[28]),
    .Q(main_basesoc_timer_reload_storage_TMR_2[29]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53413.11-53419.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[2]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[2]),
    .Q(main_basesoc_timer_reload_storage_TMR_0[2]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53413.11-53419.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[2]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[2]),
    .Q(main_basesoc_timer_reload_storage_TMR_1[2]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53413.11-53419.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[2]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[2]),
    .Q(main_basesoc_timer_reload_storage_TMR_2[2]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53609.11-53615.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[30]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[29]),
    .Q(main_basesoc_timer_reload_storage_TMR_0[30]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53609.11-53615.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[30]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[29]),
    .Q(main_basesoc_timer_reload_storage_TMR_1[30]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53609.11-53615.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[30]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[29]),
    .Q(main_basesoc_timer_reload_storage_TMR_2[30]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53616.11-53622.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[31]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[30]),
    .Q(main_basesoc_timer_reload_storage_TMR_0[31]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53616.11-53622.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[31]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[30]),
    .Q(main_basesoc_timer_reload_storage_TMR_1[31]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53616.11-53622.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[31]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[30]),
    .Q(main_basesoc_timer_reload_storage_TMR_2[31]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53420.11-53426.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[3]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[3]),
    .Q(main_basesoc_timer_reload_storage_TMR_0[3]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53420.11-53426.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[3]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[3]),
    .Q(main_basesoc_timer_reload_storage_TMR_1[3]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53420.11-53426.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[3]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[3]),
    .Q(main_basesoc_timer_reload_storage_TMR_2[3]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53427.11-53433.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[4]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[4]),
    .Q(main_basesoc_timer_reload_storage_TMR_0[4]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53427.11-53433.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[4]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[4]),
    .Q(main_basesoc_timer_reload_storage_TMR_1[4]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53427.11-53433.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[4]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[4]),
    .Q(main_basesoc_timer_reload_storage_TMR_2[4]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53434.11-53440.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[5]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[5]),
    .Q(main_basesoc_timer_reload_storage_TMR_0[5]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53434.11-53440.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[5]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[5]),
    .Q(main_basesoc_timer_reload_storage_TMR_1[5]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53434.11-53440.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[5]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[5]),
    .Q(main_basesoc_timer_reload_storage_TMR_2[5]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53441.11-53447.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[6]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[6]),
    .Q(main_basesoc_timer_reload_storage_TMR_0[6]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53441.11-53447.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[6]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[6]),
    .Q(main_basesoc_timer_reload_storage_TMR_1[6]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53441.11-53447.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[6]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[6]),
    .Q(main_basesoc_timer_reload_storage_TMR_2[6]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53448.11-53454.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[7]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[7]),
    .Q(main_basesoc_timer_reload_storage_TMR_0[7]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53448.11-53454.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[7]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[7]),
    .Q(main_basesoc_timer_reload_storage_TMR_1[7]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53448.11-53454.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[7]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[7]),
    .Q(main_basesoc_timer_reload_storage_TMR_2[7]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53455.11-53461.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[8]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[8]),
    .Q(main_basesoc_timer_reload_storage_TMR_0[8]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53455.11-53461.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[8]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[8]),
    .Q(main_basesoc_timer_reload_storage_TMR_1[8]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53455.11-53461.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[8]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[8]),
    .Q(main_basesoc_timer_reload_storage_TMR_2[8]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53462.11-53468.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[9]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[9]),
    .Q(main_basesoc_timer_reload_storage_TMR_0[9]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53462.11-53468.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[9]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[9]),
    .Q(main_basesoc_timer_reload_storage_TMR_1[9]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53462.11-53468.2" *)
  FD1P3IX \main_basesoc_timer_reload_storage_reg[9]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[9]),
    .Q(main_basesoc_timer_reload_storage_TMR_2[9]),
    .SP(builder_csr_bankarray_csrbank2_reload0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53392.11-53398.2" *)
  FD1P3IX main_basesoc_timer_update_value_re_reg_TMR_0 (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_timer_update_value_storage_0_sqmuxa_TMR_0),
    .Q(main_basesoc_timer_update_value_re_TMR_0),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53392.11-53398.2" *)
  FD1P3IX main_basesoc_timer_update_value_re_reg_TMR_1 (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_timer_update_value_storage_0_sqmuxa_TMR_1),
    .Q(main_basesoc_timer_update_value_re_TMR_1),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53392.11-53398.2" *)
  FD1P3IX main_basesoc_timer_update_value_re_reg_TMR_2 (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_timer_update_value_storage_0_sqmuxa_TMR_2),
    .Q(main_basesoc_timer_update_value_re_TMR_2),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53385.11-53391.2" *)
  FD1P3IX main_basesoc_timer_update_value_storage_reg_TMR_0 (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[0]),
    .Q(main_basesoc_timer_update_value_storage_TMR_0),
    .SP(builder_csr_bankarray_csrbank2_update_value0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53385.11-53391.2" *)
  FD1P3IX main_basesoc_timer_update_value_storage_reg_TMR_1 (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[0]),
    .Q(main_basesoc_timer_update_value_storage_TMR_1),
    .SP(builder_csr_bankarray_csrbank2_update_value0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53385.11-53391.2" *)
  FD1P3IX main_basesoc_timer_update_value_storage_reg_TMR_2 (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[0]),
    .Q(main_basesoc_timer_update_value_storage_TMR_2),
    .SP(builder_csr_bankarray_csrbank2_update_value0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53161.11-53167.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[0]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_timer_value_0_mod_RNO_TMR_0),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_0_0_TMR_0 ),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53161.11-53167.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[0]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_timer_value_0_mod_RNO_TMR_1),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_0_0_TMR_1 ),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53161.11-53167.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[0]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_timer_value_0_mod_RNO_TMR_2),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_0_0_TMR_2 ),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53231.11-53237.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[10]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_0 [10]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [10]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53231.11-53237.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[10]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_1 [10]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [10]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53231.11-53237.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[10]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_2 [10]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [10]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53238.11-53244.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[11]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_0 [11]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [11]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53238.11-53244.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[11]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_1 [11]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [11]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53238.11-53244.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[11]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_2 [11]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [11]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53245.11-53251.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[12]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_0 [12]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [12]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53245.11-53251.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[12]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_1 [12]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [12]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53245.11-53251.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[12]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_2 [12]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [12]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53252.11-53258.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[13]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_0 [13]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [13]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53252.11-53258.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[13]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_1 [13]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [13]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53252.11-53258.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[13]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_2 [13]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [13]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53259.11-53265.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[14]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_0 [14]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [14]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53259.11-53265.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[14]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_1 [14]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [14]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53259.11-53265.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[14]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_2 [14]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [14]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53266.11-53272.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[15]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_0 [15]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [15]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53266.11-53272.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[15]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_1 [15]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [15]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53266.11-53272.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[15]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_2 [15]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [15]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53273.11-53279.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[16]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_0 [16]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [16]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53273.11-53279.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[16]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_1 [16]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [16]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53273.11-53279.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[16]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_2 [16]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [16]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53280.11-53286.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[17]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_0 [17]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [17]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53280.11-53286.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[17]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_1 [17]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [17]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53280.11-53286.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[17]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_2 [17]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [17]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53287.11-53293.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[18]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_0 [18]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [18]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53287.11-53293.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[18]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_1 [18]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [18]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53287.11-53293.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[18]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_2 [18]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [18]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53294.11-53300.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[19]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_0 [19]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [19]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53294.11-53300.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[19]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_1 [19]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [19]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53294.11-53300.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[19]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_2 [19]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [19]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53168.11-53174.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[1]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_0 [1]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [1]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53168.11-53174.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[1]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_1 [1]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [1]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53168.11-53174.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[1]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_2 [1]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [1]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53301.11-53307.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[20]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_0 [20]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [20]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53301.11-53307.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[20]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_1 [20]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [20]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53301.11-53307.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[20]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_2 [20]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [20]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53308.11-53314.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[21]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_0 [21]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [21]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53308.11-53314.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[21]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_1 [21]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [21]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53308.11-53314.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[21]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_2 [21]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [21]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53315.11-53321.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[22]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_0 [22]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [22]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53315.11-53321.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[22]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_1 [22]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [22]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53315.11-53321.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[22]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_2 [22]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [22]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53322.11-53328.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[23]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_0 [23]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [23]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53322.11-53328.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[23]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_1 [23]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [23]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53322.11-53328.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[23]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_2 [23]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [23]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53329.11-53335.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[24]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_0 [24]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [24]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53329.11-53335.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[24]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_1 [24]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [24]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53329.11-53335.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[24]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_2 [24]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [24]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53336.11-53342.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[25]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_0 [25]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [25]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53336.11-53342.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[25]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_1 [25]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [25]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53336.11-53342.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[25]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_2 [25]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [25]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53343.11-53349.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[26]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_0 [26]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [26]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53343.11-53349.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[26]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_1 [26]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [26]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53343.11-53349.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[26]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_2 [26]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [26]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53350.11-53356.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[27]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_0 [27]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [27]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53350.11-53356.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[27]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_1 [27]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [27]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53350.11-53356.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[27]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_2 [27]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [27]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53357.11-53363.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[28]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_0 [28]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [28]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53357.11-53363.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[28]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_1 [28]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [28]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53357.11-53363.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[28]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_2 [28]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [28]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53364.11-53370.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[29]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_0 [29]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [29]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53364.11-53370.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[29]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_1 [29]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [29]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53364.11-53370.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[29]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_2 [29]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [29]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53175.11-53181.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[2]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_0 [2]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [2]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53175.11-53181.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[2]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_1 [2]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [2]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53175.11-53181.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[2]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_2 [2]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [2]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53371.11-53377.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[30]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_0 [30]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [30]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53371.11-53377.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[30]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_1 [30]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [30]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53371.11-53377.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[30]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_2 [30]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [30]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53378.11-53384.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[31]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_0 [31]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [31]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53378.11-53384.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[31]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_1 [31]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [31]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53378.11-53384.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[31]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_2 [31]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [31]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53182.11-53188.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[3]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_0 [3]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [3]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53182.11-53188.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[3]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_1 [3]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [3]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53182.11-53188.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[3]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_2 [3]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [3]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53189.11-53195.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[4]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_0 [4]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [4]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53189.11-53195.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[4]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_1 [4]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [4]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53189.11-53195.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[4]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_2 [4]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [4]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53196.11-53202.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[5]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_0 [5]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [5]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53196.11-53202.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[5]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_1 [5]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [5]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53196.11-53202.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[5]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_2 [5]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [5]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53203.11-53209.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[6]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_0 [6]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [6]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53203.11-53209.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[6]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_1 [6]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [6]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53203.11-53209.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[6]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_2 [6]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [6]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53210.11-53216.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[7]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_0 [7]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [7]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53210.11-53216.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[7]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_1 [7]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [7]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53210.11-53216.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[7]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_2 [7]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [7]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53217.11-53223.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[8]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_0 [8]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [8]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53217.11-53223.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[8]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_1 [8]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [8]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53217.11-53223.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[8]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_2 [8]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [8]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53224.11-53230.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[9]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_0 [9]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [9]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53224.11-53230.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[9]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_1 [9]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [9]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53224.11-53230.2" *)
  FD1P3IX \main_basesoc_timer_value_0_mod[9]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_TMR_2 [9]),
    .Q(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [9]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55621.8-55627.2" *)
  LUT4 \main_basesoc_timer_value_0_mod_RNO_cZ[0]_TMR_0  (
    .A(N_792_TMR_0),
    .B(sys_rst_TMR_0),
    .C(dsp_join_kb_TMR_0[0]),
    .D(main_basesoc_timer_en_storage_TMR_0),
    .Z(main_basesoc_timer_value_0_mod_RNO_TMR_0)
  );
  defparam \main_basesoc_timer_value_0_mod_RNO_cZ[0]_TMR_0 .INIT = "0x2230";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55621.8-55627.2" *)
  LUT4 \main_basesoc_timer_value_0_mod_RNO_cZ[0]_TMR_1  (
    .A(N_792_TMR_1),
    .B(sys_rst_TMR_1),
    .C(dsp_join_kb_TMR_1[0]),
    .D(main_basesoc_timer_en_storage_TMR_1),
    .Z(main_basesoc_timer_value_0_mod_RNO_TMR_1)
  );
  defparam \main_basesoc_timer_value_0_mod_RNO_cZ[0]_TMR_1 .INIT = "0x2230";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55621.8-55627.2" *)
  LUT4 \main_basesoc_timer_value_0_mod_RNO_cZ[0]_TMR_2  (
    .A(N_792_TMR_2),
    .B(sys_rst_TMR_2),
    .C(dsp_join_kb_TMR_2[0]),
    .D(main_basesoc_timer_en_storage_TMR_2),
    .Z(main_basesoc_timer_value_0_mod_RNO_TMR_2)
  );
  defparam \main_basesoc_timer_value_0_mod_RNO_cZ[0]_TMR_2 .INIT = "0x2230";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52937.11-52943.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[0]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_0_0_TMR_0 ),
    .Q(main_basesoc_timer_value_status_TMR_0[0]),
    .SP(main_basesoc_timer_update_value_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52937.11-52943.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[0]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_0_0_TMR_1 ),
    .Q(main_basesoc_timer_value_status_TMR_1[0]),
    .SP(main_basesoc_timer_update_value_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52937.11-52943.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[0]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_0_0_TMR_2 ),
    .Q(main_basesoc_timer_value_status_TMR_2[0]),
    .SP(main_basesoc_timer_update_value_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53007.11-53013.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[10]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [10]),
    .Q(main_basesoc_timer_value_status_TMR_0[10]),
    .SP(main_basesoc_timer_update_value_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53007.11-53013.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[10]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [10]),
    .Q(main_basesoc_timer_value_status_TMR_1[10]),
    .SP(main_basesoc_timer_update_value_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53007.11-53013.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[10]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [10]),
    .Q(main_basesoc_timer_value_status_TMR_2[10]),
    .SP(main_basesoc_timer_update_value_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53014.11-53020.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[11]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [11]),
    .Q(main_basesoc_timer_value_status_TMR_0[11]),
    .SP(main_basesoc_timer_update_value_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53014.11-53020.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[11]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [11]),
    .Q(main_basesoc_timer_value_status_TMR_1[11]),
    .SP(main_basesoc_timer_update_value_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53014.11-53020.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[11]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [11]),
    .Q(main_basesoc_timer_value_status_TMR_2[11]),
    .SP(main_basesoc_timer_update_value_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53021.11-53027.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[12]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [12]),
    .Q(main_basesoc_timer_value_status_TMR_0[12]),
    .SP(main_basesoc_timer_update_value_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53021.11-53027.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[12]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [12]),
    .Q(main_basesoc_timer_value_status_TMR_1[12]),
    .SP(main_basesoc_timer_update_value_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53021.11-53027.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[12]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [12]),
    .Q(main_basesoc_timer_value_status_TMR_2[12]),
    .SP(main_basesoc_timer_update_value_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53028.11-53034.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[13]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [13]),
    .Q(main_basesoc_timer_value_status_TMR_0[13]),
    .SP(main_basesoc_timer_update_value_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53028.11-53034.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[13]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [13]),
    .Q(main_basesoc_timer_value_status_TMR_1[13]),
    .SP(main_basesoc_timer_update_value_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53028.11-53034.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[13]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [13]),
    .Q(main_basesoc_timer_value_status_TMR_2[13]),
    .SP(main_basesoc_timer_update_value_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53035.11-53041.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[14]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [14]),
    .Q(main_basesoc_timer_value_status_TMR_0[14]),
    .SP(main_basesoc_timer_update_value_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53035.11-53041.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[14]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [14]),
    .Q(main_basesoc_timer_value_status_TMR_1[14]),
    .SP(main_basesoc_timer_update_value_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53035.11-53041.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[14]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [14]),
    .Q(main_basesoc_timer_value_status_TMR_2[14]),
    .SP(main_basesoc_timer_update_value_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53042.11-53048.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[15]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [15]),
    .Q(main_basesoc_timer_value_status_TMR_0[15]),
    .SP(main_basesoc_timer_update_value_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53042.11-53048.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[15]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [15]),
    .Q(main_basesoc_timer_value_status_TMR_1[15]),
    .SP(main_basesoc_timer_update_value_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53042.11-53048.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[15]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [15]),
    .Q(main_basesoc_timer_value_status_TMR_2[15]),
    .SP(main_basesoc_timer_update_value_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53049.11-53055.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[16]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [16]),
    .Q(main_basesoc_timer_value_status_TMR_0[16]),
    .SP(main_basesoc_timer_update_value_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53049.11-53055.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[16]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [16]),
    .Q(main_basesoc_timer_value_status_TMR_1[16]),
    .SP(main_basesoc_timer_update_value_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53049.11-53055.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[16]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [16]),
    .Q(main_basesoc_timer_value_status_TMR_2[16]),
    .SP(main_basesoc_timer_update_value_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53056.11-53062.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[17]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [17]),
    .Q(main_basesoc_timer_value_status_TMR_0[17]),
    .SP(main_basesoc_timer_update_value_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53056.11-53062.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[17]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [17]),
    .Q(main_basesoc_timer_value_status_TMR_1[17]),
    .SP(main_basesoc_timer_update_value_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53056.11-53062.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[17]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [17]),
    .Q(main_basesoc_timer_value_status_TMR_2[17]),
    .SP(main_basesoc_timer_update_value_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53063.11-53069.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[18]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [18]),
    .Q(main_basesoc_timer_value_status_TMR_0[18]),
    .SP(main_basesoc_timer_update_value_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53063.11-53069.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[18]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [18]),
    .Q(main_basesoc_timer_value_status_TMR_1[18]),
    .SP(main_basesoc_timer_update_value_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53063.11-53069.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[18]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [18]),
    .Q(main_basesoc_timer_value_status_TMR_2[18]),
    .SP(main_basesoc_timer_update_value_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53070.11-53076.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[19]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [19]),
    .Q(main_basesoc_timer_value_status_TMR_0[19]),
    .SP(main_basesoc_timer_update_value_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53070.11-53076.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[19]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [19]),
    .Q(main_basesoc_timer_value_status_TMR_1[19]),
    .SP(main_basesoc_timer_update_value_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53070.11-53076.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[19]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [19]),
    .Q(main_basesoc_timer_value_status_TMR_2[19]),
    .SP(main_basesoc_timer_update_value_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52944.11-52950.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[1]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [1]),
    .Q(main_basesoc_timer_value_status_TMR_0[1]),
    .SP(main_basesoc_timer_update_value_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52944.11-52950.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[1]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [1]),
    .Q(main_basesoc_timer_value_status_TMR_1[1]),
    .SP(main_basesoc_timer_update_value_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52944.11-52950.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[1]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [1]),
    .Q(main_basesoc_timer_value_status_TMR_2[1]),
    .SP(main_basesoc_timer_update_value_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53077.11-53083.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[20]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [20]),
    .Q(main_basesoc_timer_value_status_TMR_0[20]),
    .SP(main_basesoc_timer_update_value_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53077.11-53083.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[20]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [20]),
    .Q(main_basesoc_timer_value_status_TMR_1[20]),
    .SP(main_basesoc_timer_update_value_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53077.11-53083.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[20]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [20]),
    .Q(main_basesoc_timer_value_status_TMR_2[20]),
    .SP(main_basesoc_timer_update_value_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53084.11-53090.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[21]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [21]),
    .Q(main_basesoc_timer_value_status_TMR_0[21]),
    .SP(main_basesoc_timer_update_value_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53084.11-53090.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[21]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [21]),
    .Q(main_basesoc_timer_value_status_TMR_1[21]),
    .SP(main_basesoc_timer_update_value_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53084.11-53090.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[21]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [21]),
    .Q(main_basesoc_timer_value_status_TMR_2[21]),
    .SP(main_basesoc_timer_update_value_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53091.11-53097.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[22]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [22]),
    .Q(main_basesoc_timer_value_status_TMR_0[22]),
    .SP(main_basesoc_timer_update_value_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53091.11-53097.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[22]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [22]),
    .Q(main_basesoc_timer_value_status_TMR_1[22]),
    .SP(main_basesoc_timer_update_value_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53091.11-53097.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[22]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [22]),
    .Q(main_basesoc_timer_value_status_TMR_2[22]),
    .SP(main_basesoc_timer_update_value_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53098.11-53104.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[23]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [23]),
    .Q(main_basesoc_timer_value_status_TMR_0[23]),
    .SP(main_basesoc_timer_update_value_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53098.11-53104.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[23]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [23]),
    .Q(main_basesoc_timer_value_status_TMR_1[23]),
    .SP(main_basesoc_timer_update_value_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53098.11-53104.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[23]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [23]),
    .Q(main_basesoc_timer_value_status_TMR_2[23]),
    .SP(main_basesoc_timer_update_value_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53105.11-53111.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[24]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [24]),
    .Q(main_basesoc_timer_value_status_TMR_0[24]),
    .SP(main_basesoc_timer_update_value_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53105.11-53111.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[24]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [24]),
    .Q(main_basesoc_timer_value_status_TMR_1[24]),
    .SP(main_basesoc_timer_update_value_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53105.11-53111.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[24]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [24]),
    .Q(main_basesoc_timer_value_status_TMR_2[24]),
    .SP(main_basesoc_timer_update_value_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53112.11-53118.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[25]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [25]),
    .Q(main_basesoc_timer_value_status_TMR_0[25]),
    .SP(main_basesoc_timer_update_value_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53112.11-53118.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[25]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [25]),
    .Q(main_basesoc_timer_value_status_TMR_1[25]),
    .SP(main_basesoc_timer_update_value_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53112.11-53118.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[25]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [25]),
    .Q(main_basesoc_timer_value_status_TMR_2[25]),
    .SP(main_basesoc_timer_update_value_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53119.11-53125.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[26]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [26]),
    .Q(main_basesoc_timer_value_status_TMR_0[26]),
    .SP(main_basesoc_timer_update_value_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53119.11-53125.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[26]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [26]),
    .Q(main_basesoc_timer_value_status_TMR_1[26]),
    .SP(main_basesoc_timer_update_value_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53119.11-53125.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[26]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [26]),
    .Q(main_basesoc_timer_value_status_TMR_2[26]),
    .SP(main_basesoc_timer_update_value_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53126.11-53132.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[27]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [27]),
    .Q(main_basesoc_timer_value_status_TMR_0[27]),
    .SP(main_basesoc_timer_update_value_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53126.11-53132.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[27]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [27]),
    .Q(main_basesoc_timer_value_status_TMR_1[27]),
    .SP(main_basesoc_timer_update_value_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53126.11-53132.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[27]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [27]),
    .Q(main_basesoc_timer_value_status_TMR_2[27]),
    .SP(main_basesoc_timer_update_value_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53133.11-53139.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[28]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [28]),
    .Q(main_basesoc_timer_value_status_TMR_0[28]),
    .SP(main_basesoc_timer_update_value_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53133.11-53139.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[28]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [28]),
    .Q(main_basesoc_timer_value_status_TMR_1[28]),
    .SP(main_basesoc_timer_update_value_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53133.11-53139.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[28]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [28]),
    .Q(main_basesoc_timer_value_status_TMR_2[28]),
    .SP(main_basesoc_timer_update_value_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53140.11-53146.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[29]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [29]),
    .Q(main_basesoc_timer_value_status_TMR_0[29]),
    .SP(main_basesoc_timer_update_value_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53140.11-53146.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[29]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [29]),
    .Q(main_basesoc_timer_value_status_TMR_1[29]),
    .SP(main_basesoc_timer_update_value_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53140.11-53146.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[29]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [29]),
    .Q(main_basesoc_timer_value_status_TMR_2[29]),
    .SP(main_basesoc_timer_update_value_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52951.11-52957.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[2]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [2]),
    .Q(main_basesoc_timer_value_status_TMR_0[2]),
    .SP(main_basesoc_timer_update_value_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52951.11-52957.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[2]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [2]),
    .Q(main_basesoc_timer_value_status_TMR_1[2]),
    .SP(main_basesoc_timer_update_value_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52951.11-52957.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[2]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [2]),
    .Q(main_basesoc_timer_value_status_TMR_2[2]),
    .SP(main_basesoc_timer_update_value_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53147.11-53153.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[30]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [30]),
    .Q(main_basesoc_timer_value_status_TMR_0[30]),
    .SP(main_basesoc_timer_update_value_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53147.11-53153.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[30]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [30]),
    .Q(main_basesoc_timer_value_status_TMR_1[30]),
    .SP(main_basesoc_timer_update_value_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53147.11-53153.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[30]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [30]),
    .Q(main_basesoc_timer_value_status_TMR_2[30]),
    .SP(main_basesoc_timer_update_value_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53154.11-53160.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[31]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [31]),
    .Q(main_basesoc_timer_value_status_TMR_0[31]),
    .SP(main_basesoc_timer_update_value_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53154.11-53160.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[31]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [31]),
    .Q(main_basesoc_timer_value_status_TMR_1[31]),
    .SP(main_basesoc_timer_update_value_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53154.11-53160.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[31]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [31]),
    .Q(main_basesoc_timer_value_status_TMR_2[31]),
    .SP(main_basesoc_timer_update_value_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52958.11-52964.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[3]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [3]),
    .Q(main_basesoc_timer_value_status_TMR_0[3]),
    .SP(main_basesoc_timer_update_value_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52958.11-52964.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[3]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [3]),
    .Q(main_basesoc_timer_value_status_TMR_1[3]),
    .SP(main_basesoc_timer_update_value_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52958.11-52964.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[3]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [3]),
    .Q(main_basesoc_timer_value_status_TMR_2[3]),
    .SP(main_basesoc_timer_update_value_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52965.11-52971.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[4]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [4]),
    .Q(main_basesoc_timer_value_status_TMR_0[4]),
    .SP(main_basesoc_timer_update_value_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52965.11-52971.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[4]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [4]),
    .Q(main_basesoc_timer_value_status_TMR_1[4]),
    .SP(main_basesoc_timer_update_value_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52965.11-52971.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[4]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [4]),
    .Q(main_basesoc_timer_value_status_TMR_2[4]),
    .SP(main_basesoc_timer_update_value_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52972.11-52978.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[5]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [5]),
    .Q(main_basesoc_timer_value_status_TMR_0[5]),
    .SP(main_basesoc_timer_update_value_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52972.11-52978.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[5]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [5]),
    .Q(main_basesoc_timer_value_status_TMR_1[5]),
    .SP(main_basesoc_timer_update_value_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52972.11-52978.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[5]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [5]),
    .Q(main_basesoc_timer_value_status_TMR_2[5]),
    .SP(main_basesoc_timer_update_value_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52979.11-52985.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[6]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [6]),
    .Q(main_basesoc_timer_value_status_TMR_0[6]),
    .SP(main_basesoc_timer_update_value_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52979.11-52985.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[6]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [6]),
    .Q(main_basesoc_timer_value_status_TMR_1[6]),
    .SP(main_basesoc_timer_update_value_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52979.11-52985.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[6]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [6]),
    .Q(main_basesoc_timer_value_status_TMR_2[6]),
    .SP(main_basesoc_timer_update_value_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52986.11-52992.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[7]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [7]),
    .Q(main_basesoc_timer_value_status_TMR_0[7]),
    .SP(main_basesoc_timer_update_value_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52986.11-52992.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[7]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [7]),
    .Q(main_basesoc_timer_value_status_TMR_1[7]),
    .SP(main_basesoc_timer_update_value_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52986.11-52992.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[7]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [7]),
    .Q(main_basesoc_timer_value_status_TMR_2[7]),
    .SP(main_basesoc_timer_update_value_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52993.11-52999.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[8]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [8]),
    .Q(main_basesoc_timer_value_status_TMR_0[8]),
    .SP(main_basesoc_timer_update_value_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52993.11-52999.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[8]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [8]),
    .Q(main_basesoc_timer_value_status_TMR_1[8]),
    .SP(main_basesoc_timer_update_value_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52993.11-52999.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[8]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [8]),
    .Q(main_basesoc_timer_value_status_TMR_2[8]),
    .SP(main_basesoc_timer_update_value_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53000.11-53006.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[9]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_0 [9]),
    .Q(main_basesoc_timer_value_status_TMR_0[9]),
    .SP(main_basesoc_timer_update_value_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53000.11-53006.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[9]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_1 [9]),
    .Q(main_basesoc_timer_value_status_TMR_1[9]),
    .SP(main_basesoc_timer_update_value_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:53000.11-53006.2" *)
  FD1P3IX \main_basesoc_timer_value_status_reg[9]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\VexRiscv.IBusCachedPlugin_cache.main_basesoc_timer_value_7_1_TMR_2 [9]),
    .Q(main_basesoc_timer_value_status_TMR_2[9]),
    .SP(main_basesoc_timer_update_value_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52930.11-52936.2" *)
  FD1P3IX main_basesoc_timer_zero_pending_reg_TMR_0 (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(N_136_TMR_0),
    .Q(main_basesoc_timer_zero_pending_TMR_0),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52930.11-52936.2" *)
  FD1P3IX main_basesoc_timer_zero_pending_reg_TMR_1 (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(N_136_TMR_1),
    .Q(main_basesoc_timer_zero_pending_TMR_1),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52930.11-52936.2" *)
  FD1P3IX main_basesoc_timer_zero_pending_reg_TMR_2 (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(N_136_TMR_2),
    .Q(main_basesoc_timer_zero_pending_TMR_2),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52923.11-52929.2" *)
  FD1P3IX main_basesoc_timer_zero_trigger_d_reg_TMR_0 (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(main_basesoc_timer_zero_trigger_TMR_0),
    .Q(main_basesoc_timer_zero_trigger_d_TMR_0),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52923.11-52929.2" *)
  FD1P3IX main_basesoc_timer_zero_trigger_d_reg_TMR_1 (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(main_basesoc_timer_zero_trigger_TMR_1),
    .Q(main_basesoc_timer_zero_trigger_d_TMR_1),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52923.11-52929.2" *)
  FD1P3IX main_basesoc_timer_zero_trigger_d_reg_TMR_2 (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(main_basesoc_timer_zero_trigger_TMR_2),
    .Q(main_basesoc_timer_zero_trigger_d_TMR_2),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52895.11-52901.2" *)
  FD1P3IX \main_basesoc_tx_count[0]_TMR_0  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_0),
    .CK(sys_clk),
    .D(\main_basesoc_tx_count_0_.fb_TMR_0 ),
    .Q(CO0_0_TMR_0),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52895.11-52901.2" *)
  FD1P3IX \main_basesoc_tx_count[0]_TMR_1  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_1),
    .CK(sys_clk),
    .D(\main_basesoc_tx_count_0_.fb_TMR_1 ),
    .Q(CO0_0_TMR_1),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52895.11-52901.2" *)
  FD1P3IX \main_basesoc_tx_count[0]_TMR_2  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_2),
    .CK(sys_clk),
    .D(\main_basesoc_tx_count_0_.fb_TMR_2 ),
    .Q(CO0_0_TMR_2),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51398.8-51404.2" *)
  LUT4 \main_basesoc_tx_count_0_.fb_cZ_TMR_0  (
    .A(CO0_0_TMR_0),
    .B(main_basesoc_tx_tick_TMR_0),
    .C(builder_basesoc_rs232phytx_state_TMR_0),
    .D(GND_0),
    .Z(\main_basesoc_tx_count_0_.fb_TMR_0 )
  );
  defparam \main_basesoc_tx_count_0_.fb_cZ_TMR_0 .INIT = "0x6565";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51398.8-51404.2" *)
  LUT4 \main_basesoc_tx_count_0_.fb_cZ_TMR_1  (
    .A(CO0_0_TMR_1),
    .B(main_basesoc_tx_tick_TMR_1),
    .C(builder_basesoc_rs232phytx_state_TMR_1),
    .D(GND_0),
    .Z(\main_basesoc_tx_count_0_.fb_TMR_1 )
  );
  defparam \main_basesoc_tx_count_0_.fb_cZ_TMR_1 .INIT = "0x6565";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51398.8-51404.2" *)
  LUT4 \main_basesoc_tx_count_0_.fb_cZ_TMR_2  (
    .A(CO0_0_TMR_2),
    .B(main_basesoc_tx_tick_TMR_2),
    .C(builder_basesoc_rs232phytx_state_TMR_2),
    .D(GND_0),
    .Z(\main_basesoc_tx_count_0_.fb_TMR_2 )
  );
  defparam \main_basesoc_tx_count_0_.fb_cZ_TMR_2 .INIT = "0x6565";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52902.11-52908.2" *)
  FD1P3IX \main_basesoc_tx_count_reg[1]_TMR_0  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_0),
    .CK(sys_clk),
    .D(main_basesoc_tx_count_rs232phytx_next_value0_TMR_0[1]),
    .Q(main_basesoc_tx_count_TMR_0[1]),
    .SP(main_basesoc_serial_tx_rs232phytx_next_value1_1_sqmuxa_i_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52902.11-52908.2" *)
  FD1P3IX \main_basesoc_tx_count_reg[1]_TMR_1  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_1),
    .CK(sys_clk),
    .D(main_basesoc_tx_count_rs232phytx_next_value0_TMR_1[1]),
    .Q(main_basesoc_tx_count_TMR_1[1]),
    .SP(main_basesoc_serial_tx_rs232phytx_next_value1_1_sqmuxa_i_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52902.11-52908.2" *)
  FD1P3IX \main_basesoc_tx_count_reg[1]_TMR_2  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_2),
    .CK(sys_clk),
    .D(main_basesoc_tx_count_rs232phytx_next_value0_TMR_2[1]),
    .Q(main_basesoc_tx_count_TMR_2[1]),
    .SP(main_basesoc_serial_tx_rs232phytx_next_value1_1_sqmuxa_i_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52909.11-52915.2" *)
  FD1P3IX \main_basesoc_tx_count_reg[2]_TMR_0  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_0),
    .CK(sys_clk),
    .D(main_basesoc_tx_count_rs232phytx_next_value0_TMR_0[2]),
    .Q(main_basesoc_tx_count_TMR_0[2]),
    .SP(main_basesoc_serial_tx_rs232phytx_next_value1_1_sqmuxa_i_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52909.11-52915.2" *)
  FD1P3IX \main_basesoc_tx_count_reg[2]_TMR_1  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_1),
    .CK(sys_clk),
    .D(main_basesoc_tx_count_rs232phytx_next_value0_TMR_1[2]),
    .Q(main_basesoc_tx_count_TMR_1[2]),
    .SP(main_basesoc_serial_tx_rs232phytx_next_value1_1_sqmuxa_i_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52909.11-52915.2" *)
  FD1P3IX \main_basesoc_tx_count_reg[2]_TMR_2  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_2),
    .CK(sys_clk),
    .D(main_basesoc_tx_count_rs232phytx_next_value0_TMR_2[2]),
    .Q(main_basesoc_tx_count_TMR_2[2]),
    .SP(main_basesoc_serial_tx_rs232phytx_next_value1_1_sqmuxa_i_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52916.11-52922.2" *)
  FD1P3IX \main_basesoc_tx_count_reg[3]_TMR_0  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_0),
    .CK(sys_clk),
    .D(main_basesoc_tx_count_rs232phytx_next_value0_TMR_0[3]),
    .Q(main_basesoc_tx_count_TMR_0[3]),
    .SP(main_basesoc_serial_tx_rs232phytx_next_value1_1_sqmuxa_i_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52916.11-52922.2" *)
  FD1P3IX \main_basesoc_tx_count_reg[3]_TMR_1  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_1),
    .CK(sys_clk),
    .D(main_basesoc_tx_count_rs232phytx_next_value0_TMR_1[3]),
    .Q(main_basesoc_tx_count_TMR_1[3]),
    .SP(main_basesoc_serial_tx_rs232phytx_next_value1_1_sqmuxa_i_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52916.11-52922.2" *)
  FD1P3IX \main_basesoc_tx_count_reg[3]_TMR_2  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_2),
    .CK(sys_clk),
    .D(main_basesoc_tx_count_rs232phytx_next_value0_TMR_2[3]),
    .Q(main_basesoc_tx_count_TMR_2[3]),
    .SP(main_basesoc_serial_tx_rs232phytx_next_value1_1_sqmuxa_i_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52839.11-52845.2" *)
  FD1P3IX \main_basesoc_tx_data_reg[0]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_tx_data_rs232phytx_next_value2_TMR_0[0]),
    .Q(main_basesoc_tx_data_TMR_0[0]),
    .SP(main_basesoc_tx_data_rs232phytx_next_value_ce2_1_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52839.11-52845.2" *)
  FD1P3IX \main_basesoc_tx_data_reg[0]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_tx_data_rs232phytx_next_value2_TMR_1[0]),
    .Q(main_basesoc_tx_data_TMR_1[0]),
    .SP(main_basesoc_tx_data_rs232phytx_next_value_ce2_1_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52839.11-52845.2" *)
  FD1P3IX \main_basesoc_tx_data_reg[0]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_tx_data_rs232phytx_next_value2_TMR_2[0]),
    .Q(main_basesoc_tx_data_TMR_2[0]),
    .SP(main_basesoc_tx_data_rs232phytx_next_value_ce2_1_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52846.11-52852.2" *)
  FD1P3IX \main_basesoc_tx_data_reg[1]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_tx_data_rs232phytx_next_value2_TMR_0[1]),
    .Q(main_basesoc_tx_data_TMR_0[1]),
    .SP(main_basesoc_tx_data_rs232phytx_next_value_ce2_1_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52846.11-52852.2" *)
  FD1P3IX \main_basesoc_tx_data_reg[1]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_tx_data_rs232phytx_next_value2_TMR_1[1]),
    .Q(main_basesoc_tx_data_TMR_1[1]),
    .SP(main_basesoc_tx_data_rs232phytx_next_value_ce2_1_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52846.11-52852.2" *)
  FD1P3IX \main_basesoc_tx_data_reg[1]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_tx_data_rs232phytx_next_value2_TMR_2[1]),
    .Q(main_basesoc_tx_data_TMR_2[1]),
    .SP(main_basesoc_tx_data_rs232phytx_next_value_ce2_1_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52853.11-52859.2" *)
  FD1P3IX \main_basesoc_tx_data_reg[2]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_tx_data_rs232phytx_next_value2_TMR_0[2]),
    .Q(main_basesoc_tx_data_TMR_0[2]),
    .SP(main_basesoc_tx_data_rs232phytx_next_value_ce2_1_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52853.11-52859.2" *)
  FD1P3IX \main_basesoc_tx_data_reg[2]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_tx_data_rs232phytx_next_value2_TMR_1[2]),
    .Q(main_basesoc_tx_data_TMR_1[2]),
    .SP(main_basesoc_tx_data_rs232phytx_next_value_ce2_1_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52853.11-52859.2" *)
  FD1P3IX \main_basesoc_tx_data_reg[2]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_tx_data_rs232phytx_next_value2_TMR_2[2]),
    .Q(main_basesoc_tx_data_TMR_2[2]),
    .SP(main_basesoc_tx_data_rs232phytx_next_value_ce2_1_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52860.11-52866.2" *)
  FD1P3IX \main_basesoc_tx_data_reg[3]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_tx_data_rs232phytx_next_value2_TMR_0[3]),
    .Q(main_basesoc_tx_data_TMR_0[3]),
    .SP(main_basesoc_tx_data_rs232phytx_next_value_ce2_1_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52860.11-52866.2" *)
  FD1P3IX \main_basesoc_tx_data_reg[3]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_tx_data_rs232phytx_next_value2_TMR_1[3]),
    .Q(main_basesoc_tx_data_TMR_1[3]),
    .SP(main_basesoc_tx_data_rs232phytx_next_value_ce2_1_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52860.11-52866.2" *)
  FD1P3IX \main_basesoc_tx_data_reg[3]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_tx_data_rs232phytx_next_value2_TMR_2[3]),
    .Q(main_basesoc_tx_data_TMR_2[3]),
    .SP(main_basesoc_tx_data_rs232phytx_next_value_ce2_1_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52867.11-52873.2" *)
  FD1P3IX \main_basesoc_tx_data_reg[4]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_tx_data_rs232phytx_next_value2_TMR_0[4]),
    .Q(main_basesoc_tx_data_TMR_0[4]),
    .SP(main_basesoc_tx_data_rs232phytx_next_value_ce2_1_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52867.11-52873.2" *)
  FD1P3IX \main_basesoc_tx_data_reg[4]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_tx_data_rs232phytx_next_value2_TMR_1[4]),
    .Q(main_basesoc_tx_data_TMR_1[4]),
    .SP(main_basesoc_tx_data_rs232phytx_next_value_ce2_1_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52867.11-52873.2" *)
  FD1P3IX \main_basesoc_tx_data_reg[4]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_tx_data_rs232phytx_next_value2_TMR_2[4]),
    .Q(main_basesoc_tx_data_TMR_2[4]),
    .SP(main_basesoc_tx_data_rs232phytx_next_value_ce2_1_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52874.11-52880.2" *)
  FD1P3IX \main_basesoc_tx_data_reg[5]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_tx_data_rs232phytx_next_value2_TMR_0[5]),
    .Q(main_basesoc_tx_data_TMR_0[5]),
    .SP(main_basesoc_tx_data_rs232phytx_next_value_ce2_1_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52874.11-52880.2" *)
  FD1P3IX \main_basesoc_tx_data_reg[5]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_tx_data_rs232phytx_next_value2_TMR_1[5]),
    .Q(main_basesoc_tx_data_TMR_1[5]),
    .SP(main_basesoc_tx_data_rs232phytx_next_value_ce2_1_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52874.11-52880.2" *)
  FD1P3IX \main_basesoc_tx_data_reg[5]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_tx_data_rs232phytx_next_value2_TMR_2[5]),
    .Q(main_basesoc_tx_data_TMR_2[5]),
    .SP(main_basesoc_tx_data_rs232phytx_next_value_ce2_1_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52881.11-52887.2" *)
  FD1P3IX \main_basesoc_tx_data_reg[6]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_tx_data_rs232phytx_next_value2_TMR_0[6]),
    .Q(main_basesoc_tx_data_TMR_0[6]),
    .SP(main_basesoc_tx_data_rs232phytx_next_value_ce2_1_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52881.11-52887.2" *)
  FD1P3IX \main_basesoc_tx_data_reg[6]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_tx_data_rs232phytx_next_value2_TMR_1[6]),
    .Q(main_basesoc_tx_data_TMR_1[6]),
    .SP(main_basesoc_tx_data_rs232phytx_next_value_ce2_1_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52881.11-52887.2" *)
  FD1P3IX \main_basesoc_tx_data_reg[6]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_tx_data_rs232phytx_next_value2_TMR_2[6]),
    .Q(main_basesoc_tx_data_TMR_2[6]),
    .SP(main_basesoc_tx_data_rs232phytx_next_value_ce2_1_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52888.11-52894.2" *)
  FD1P3IX \main_basesoc_tx_data_reg[7]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_tx_data_rs232phytx_next_value2_TMR_0[7]),
    .Q(main_basesoc_tx_data_TMR_0[7]),
    .SP(main_basesoc_tx_data_rs232phytx_next_value_ce2_1_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52888.11-52894.2" *)
  FD1P3IX \main_basesoc_tx_data_reg[7]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_tx_data_rs232phytx_next_value2_TMR_1[7]),
    .Q(main_basesoc_tx_data_TMR_1[7]),
    .SP(main_basesoc_tx_data_rs232phytx_next_value_ce2_1_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52888.11-52894.2" *)
  FD1P3IX \main_basesoc_tx_data_reg[7]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_tx_data_rs232phytx_next_value2_TMR_2[7]),
    .Q(main_basesoc_tx_data_TMR_2[7]),
    .SP(main_basesoc_tx_data_rs232phytx_next_value_ce2_1_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52685.11-52691.2" *)
  FD1P3IX \main_basesoc_tx_phase[10]_TMR_0  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_0),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_9_0_S1_TMR_0),
    .Q(dsp_join_kb_26_TMR_0[10]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52685.11-52691.2" *)
  FD1P3IX \main_basesoc_tx_phase[10]_TMR_1  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_1),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_9_0_S1_TMR_1),
    .Q(dsp_join_kb_26_TMR_1[10]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52685.11-52691.2" *)
  FD1P3IX \main_basesoc_tx_phase[10]_TMR_2  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_2),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_9_0_S1_TMR_2),
    .Q(dsp_join_kb_26_TMR_2[10]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52692.11-52698.2" *)
  FD1P3IX \main_basesoc_tx_phase[11]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(N_17833_0_TMR_0),
    .Q(dsp_join_kb_26_TMR_0[11]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52692.11-52698.2" *)
  FD1P3IX \main_basesoc_tx_phase[11]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(N_17833_0_TMR_1),
    .Q(dsp_join_kb_26_TMR_1[11]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52692.11-52698.2" *)
  FD1P3IX \main_basesoc_tx_phase[11]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(N_17833_0_TMR_2),
    .Q(dsp_join_kb_26_TMR_2[11]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52699.11-52705.2" *)
  FD1P3IX \main_basesoc_tx_phase[12]_TMR_0  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_0),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_11_0_S1_TMR_0),
    .Q(dsp_join_kb_26_TMR_0[12]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52699.11-52705.2" *)
  FD1P3IX \main_basesoc_tx_phase[12]_TMR_1  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_1),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_11_0_S1_TMR_1),
    .Q(dsp_join_kb_26_TMR_1[12]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52699.11-52705.2" *)
  FD1P3IX \main_basesoc_tx_phase[12]_TMR_2  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_2),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_11_0_S1_TMR_2),
    .Q(dsp_join_kb_26_TMR_2[12]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52706.11-52712.2" *)
  FD1P3IX \main_basesoc_tx_phase[13]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(N_17835_0_TMR_0),
    .Q(dsp_join_kb_26_TMR_0[13]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52706.11-52712.2" *)
  FD1P3IX \main_basesoc_tx_phase[13]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(N_17835_0_TMR_1),
    .Q(dsp_join_kb_26_TMR_1[13]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52706.11-52712.2" *)
  FD1P3IX \main_basesoc_tx_phase[13]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(N_17835_0_TMR_2),
    .Q(dsp_join_kb_26_TMR_2[13]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52713.11-52719.2" *)
  FD1P3IX \main_basesoc_tx_phase[14]_TMR_0  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_0),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_13_0_S1_TMR_0),
    .Q(dsp_join_kb_26_TMR_0[14]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52713.11-52719.2" *)
  FD1P3IX \main_basesoc_tx_phase[14]_TMR_1  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_1),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_13_0_S1_TMR_1),
    .Q(dsp_join_kb_26_TMR_1[14]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52713.11-52719.2" *)
  FD1P3IX \main_basesoc_tx_phase[14]_TMR_2  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_2),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_13_0_S1_TMR_2),
    .Q(dsp_join_kb_26_TMR_2[14]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52720.11-52726.2" *)
  FD1P3IX \main_basesoc_tx_phase[15]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(N_17815_0_TMR_0),
    .Q(dsp_join_kb_26_TMR_0[15]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52720.11-52726.2" *)
  FD1P3IX \main_basesoc_tx_phase[15]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(N_17815_0_TMR_1),
    .Q(dsp_join_kb_26_TMR_1[15]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52720.11-52726.2" *)
  FD1P3IX \main_basesoc_tx_phase[15]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(N_17815_0_TMR_2),
    .Q(dsp_join_kb_26_TMR_2[15]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52727.11-52733.2" *)
  FD1P3IX \main_basesoc_tx_phase[16]_TMR_0  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_0),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_15_0_S1_TMR_0),
    .Q(dsp_join_kb_26_TMR_0[16]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52727.11-52733.2" *)
  FD1P3IX \main_basesoc_tx_phase[16]_TMR_1  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_1),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_15_0_S1_TMR_1),
    .Q(dsp_join_kb_26_TMR_1[16]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52727.11-52733.2" *)
  FD1P3IX \main_basesoc_tx_phase[16]_TMR_2  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_2),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_15_0_S1_TMR_2),
    .Q(dsp_join_kb_26_TMR_2[16]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52734.11-52740.2" *)
  FD1P3IX \main_basesoc_tx_phase[17]_TMR_0  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_0),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_17_0_S0_TMR_0),
    .Q(dsp_join_kb_26_TMR_0[17]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52734.11-52740.2" *)
  FD1P3IX \main_basesoc_tx_phase[17]_TMR_1  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_1),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_17_0_S0_TMR_1),
    .Q(dsp_join_kb_26_TMR_1[17]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52734.11-52740.2" *)
  FD1P3IX \main_basesoc_tx_phase[17]_TMR_2  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_2),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_17_0_S0_TMR_2),
    .Q(dsp_join_kb_26_TMR_2[17]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52741.11-52747.2" *)
  FD1P3IX \main_basesoc_tx_phase[18]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(N_17817_0_TMR_0),
    .Q(dsp_join_kb_26_TMR_0[18]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52741.11-52747.2" *)
  FD1P3IX \main_basesoc_tx_phase[18]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(N_17817_0_TMR_1),
    .Q(dsp_join_kb_26_TMR_1[18]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52741.11-52747.2" *)
  FD1P3IX \main_basesoc_tx_phase[18]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(N_17817_0_TMR_2),
    .Q(dsp_join_kb_26_TMR_2[18]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52748.11-52754.2" *)
  FD1P3IX \main_basesoc_tx_phase[19]_TMR_0  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_0),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_19_0_S0_TMR_0),
    .Q(dsp_join_kb_26_TMR_0[19]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52748.11-52754.2" *)
  FD1P3IX \main_basesoc_tx_phase[19]_TMR_1  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_1),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_19_0_S0_TMR_1),
    .Q(dsp_join_kb_26_TMR_1[19]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52748.11-52754.2" *)
  FD1P3IX \main_basesoc_tx_phase[19]_TMR_2  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_2),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_19_0_S0_TMR_2),
    .Q(dsp_join_kb_26_TMR_2[19]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52622.11-52628.2" *)
  FD1P3IX \main_basesoc_tx_phase[1]_TMR_0  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_0),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_1_0_S0_TMR_0),
    .Q(dsp_join_kb_26_TMR_0[1]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52622.11-52628.2" *)
  FD1P3IX \main_basesoc_tx_phase[1]_TMR_1  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_1),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_1_0_S0_TMR_1),
    .Q(dsp_join_kb_26_TMR_1[1]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52622.11-52628.2" *)
  FD1P3IX \main_basesoc_tx_phase[1]_TMR_2  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_2),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_1_0_S0_TMR_2),
    .Q(dsp_join_kb_26_TMR_2[1]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52755.11-52761.2" *)
  FD1P3IX \main_basesoc_tx_phase[20]_TMR_0  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_0),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_19_0_S1_TMR_0),
    .Q(dsp_join_kb_26_TMR_0[20]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52755.11-52761.2" *)
  FD1P3IX \main_basesoc_tx_phase[20]_TMR_1  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_1),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_19_0_S1_TMR_1),
    .Q(dsp_join_kb_26_TMR_1[20]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52755.11-52761.2" *)
  FD1P3IX \main_basesoc_tx_phase[20]_TMR_2  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_2),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_19_0_S1_TMR_2),
    .Q(dsp_join_kb_26_TMR_2[20]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52762.11-52768.2" *)
  FD1P3IX \main_basesoc_tx_phase[21]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(N_17819_0_TMR_0),
    .Q(dsp_join_kb_26_TMR_0[21]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52762.11-52768.2" *)
  FD1P3IX \main_basesoc_tx_phase[21]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(N_17819_0_TMR_1),
    .Q(dsp_join_kb_26_TMR_1[21]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52762.11-52768.2" *)
  FD1P3IX \main_basesoc_tx_phase[21]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(N_17819_0_TMR_2),
    .Q(dsp_join_kb_26_TMR_2[21]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52769.11-52775.2" *)
  FD1P3IX \main_basesoc_tx_phase[22]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(N_17821_0_TMR_0),
    .Q(dsp_join_kb_26_TMR_0[22]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52769.11-52775.2" *)
  FD1P3IX \main_basesoc_tx_phase[22]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(N_17821_0_TMR_1),
    .Q(dsp_join_kb_26_TMR_1[22]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52769.11-52775.2" *)
  FD1P3IX \main_basesoc_tx_phase[22]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(N_17821_0_TMR_2),
    .Q(dsp_join_kb_26_TMR_2[22]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52776.11-52782.2" *)
  FD1P3IX \main_basesoc_tx_phase[23]_TMR_0  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_0),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_23_0_S0_TMR_0),
    .Q(dsp_join_kb_26_TMR_0[23]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52776.11-52782.2" *)
  FD1P3IX \main_basesoc_tx_phase[23]_TMR_1  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_1),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_23_0_S0_TMR_1),
    .Q(dsp_join_kb_26_TMR_1[23]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52776.11-52782.2" *)
  FD1P3IX \main_basesoc_tx_phase[23]_TMR_2  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_2),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_23_0_S0_TMR_2),
    .Q(dsp_join_kb_26_TMR_2[23]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52783.11-52789.2" *)
  FD1P3IX \main_basesoc_tx_phase[24]_TMR_0  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_0),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_23_0_S1_TMR_0),
    .Q(dsp_join_kb_26_TMR_0[24]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52783.11-52789.2" *)
  FD1P3IX \main_basesoc_tx_phase[24]_TMR_1  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_1),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_23_0_S1_TMR_1),
    .Q(dsp_join_kb_26_TMR_1[24]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52783.11-52789.2" *)
  FD1P3IX \main_basesoc_tx_phase[24]_TMR_2  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_2),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_23_0_S1_TMR_2),
    .Q(dsp_join_kb_26_TMR_2[24]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52790.11-52796.2" *)
  FD1P3IX \main_basesoc_tx_phase[25]_TMR_0  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_0),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_25_0_S0_TMR_0),
    .Q(dsp_join_kb_26_TMR_0[25]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52790.11-52796.2" *)
  FD1P3IX \main_basesoc_tx_phase[25]_TMR_1  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_1),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_25_0_S0_TMR_1),
    .Q(dsp_join_kb_26_TMR_1[25]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52790.11-52796.2" *)
  FD1P3IX \main_basesoc_tx_phase[25]_TMR_2  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_2),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_25_0_S0_TMR_2),
    .Q(dsp_join_kb_26_TMR_2[25]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52797.11-52803.2" *)
  FD1P3IX \main_basesoc_tx_phase[26]_TMR_0  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_0),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_25_0_S1_TMR_0),
    .Q(dsp_join_kb_26_TMR_0[26]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52797.11-52803.2" *)
  FD1P3IX \main_basesoc_tx_phase[26]_TMR_1  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_1),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_25_0_S1_TMR_1),
    .Q(dsp_join_kb_26_TMR_1[26]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52797.11-52803.2" *)
  FD1P3IX \main_basesoc_tx_phase[26]_TMR_2  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_2),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_25_0_S1_TMR_2),
    .Q(dsp_join_kb_26_TMR_2[26]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52804.11-52810.2" *)
  FD1P3IX \main_basesoc_tx_phase[27]_TMR_0  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_0),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_27_0_S0_TMR_0),
    .Q(dsp_join_kb_26_TMR_0[27]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52804.11-52810.2" *)
  FD1P3IX \main_basesoc_tx_phase[27]_TMR_1  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_1),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_27_0_S0_TMR_1),
    .Q(dsp_join_kb_26_TMR_1[27]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52804.11-52810.2" *)
  FD1P3IX \main_basesoc_tx_phase[27]_TMR_2  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_2),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_27_0_S0_TMR_2),
    .Q(dsp_join_kb_26_TMR_2[27]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52811.11-52817.2" *)
  FD1P3IX \main_basesoc_tx_phase[28]_TMR_0  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_0),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_27_0_S1_TMR_0),
    .Q(dsp_join_kb_26_TMR_0[28]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52811.11-52817.2" *)
  FD1P3IX \main_basesoc_tx_phase[28]_TMR_1  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_1),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_27_0_S1_TMR_1),
    .Q(dsp_join_kb_26_TMR_1[28]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52811.11-52817.2" *)
  FD1P3IX \main_basesoc_tx_phase[28]_TMR_2  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_2),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_27_0_S1_TMR_2),
    .Q(dsp_join_kb_26_TMR_2[28]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52818.11-52824.2" *)
  FD1P3IX \main_basesoc_tx_phase[29]_TMR_0  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_0),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_29_0_S0_TMR_0),
    .Q(dsp_join_kb_26_TMR_0[29]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52818.11-52824.2" *)
  FD1P3IX \main_basesoc_tx_phase[29]_TMR_1  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_1),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_29_0_S0_TMR_1),
    .Q(dsp_join_kb_26_TMR_1[29]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52818.11-52824.2" *)
  FD1P3IX \main_basesoc_tx_phase[29]_TMR_2  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_2),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_29_0_S0_TMR_2),
    .Q(dsp_join_kb_26_TMR_2[29]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52629.11-52635.2" *)
  FD1P3IX \main_basesoc_tx_phase[2]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(N_17823_0_TMR_0),
    .Q(dsp_join_kb_26_TMR_0[2]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52629.11-52635.2" *)
  FD1P3IX \main_basesoc_tx_phase[2]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(N_17823_0_TMR_1),
    .Q(dsp_join_kb_26_TMR_1[2]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52629.11-52635.2" *)
  FD1P3IX \main_basesoc_tx_phase[2]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(N_17823_0_TMR_2),
    .Q(dsp_join_kb_26_TMR_2[2]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52825.11-52831.2" *)
  FD1P3IX \main_basesoc_tx_phase[30]_TMR_0  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_0),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_29_0_S1_TMR_0),
    .Q(dsp_join_kb_26_TMR_0[30]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52825.11-52831.2" *)
  FD1P3IX \main_basesoc_tx_phase[30]_TMR_1  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_1),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_29_0_S1_TMR_1),
    .Q(dsp_join_kb_26_TMR_1[30]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52825.11-52831.2" *)
  FD1P3IX \main_basesoc_tx_phase[30]_TMR_2  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_2),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_29_0_S1_TMR_2),
    .Q(dsp_join_kb_26_TMR_2[30]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52832.11-52838.2" *)
  FD1P3IX \main_basesoc_tx_phase[31]_TMR_0  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_0),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_31_0_S0_TMR_0),
    .Q(dsp_join_kb_26_TMR_0[31]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52832.11-52838.2" *)
  FD1P3IX \main_basesoc_tx_phase[31]_TMR_1  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_1),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_31_0_S0_TMR_1),
    .Q(dsp_join_kb_26_TMR_1[31]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52832.11-52838.2" *)
  FD1P3IX \main_basesoc_tx_phase[31]_TMR_2  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_2),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_31_0_S0_TMR_2),
    .Q(dsp_join_kb_26_TMR_2[31]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52636.11-52642.2" *)
  FD1P3IX \main_basesoc_tx_phase[3]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(N_17825_0_TMR_0),
    .Q(dsp_join_kb_26_TMR_0[3]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52636.11-52642.2" *)
  FD1P3IX \main_basesoc_tx_phase[3]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(N_17825_0_TMR_1),
    .Q(dsp_join_kb_26_TMR_1[3]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52636.11-52642.2" *)
  FD1P3IX \main_basesoc_tx_phase[3]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(N_17825_0_TMR_2),
    .Q(dsp_join_kb_26_TMR_2[3]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52643.11-52649.2" *)
  FD1P3IX \main_basesoc_tx_phase[4]_TMR_0  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_0),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_3_0_S1_TMR_0),
    .Q(dsp_join_kb_26_TMR_0[4]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52643.11-52649.2" *)
  FD1P3IX \main_basesoc_tx_phase[4]_TMR_1  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_1),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_3_0_S1_TMR_1),
    .Q(dsp_join_kb_26_TMR_1[4]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52643.11-52649.2" *)
  FD1P3IX \main_basesoc_tx_phase[4]_TMR_2  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_2),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_3_0_S1_TMR_2),
    .Q(dsp_join_kb_26_TMR_2[4]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52650.11-52656.2" *)
  FD1P3IX \main_basesoc_tx_phase[5]_TMR_0  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_0),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_5_0_S0_TMR_0),
    .Q(dsp_join_kb_26_TMR_0[5]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52650.11-52656.2" *)
  FD1P3IX \main_basesoc_tx_phase[5]_TMR_1  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_1),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_5_0_S0_TMR_1),
    .Q(dsp_join_kb_26_TMR_1[5]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52650.11-52656.2" *)
  FD1P3IX \main_basesoc_tx_phase[5]_TMR_2  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_2),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_5_0_S0_TMR_2),
    .Q(dsp_join_kb_26_TMR_2[5]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52657.11-52663.2" *)
  FD1P3IX \main_basesoc_tx_phase[6]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(N_17827_0_TMR_0),
    .Q(dsp_join_kb_26_TMR_0[6]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52657.11-52663.2" *)
  FD1P3IX \main_basesoc_tx_phase[6]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(N_17827_0_TMR_1),
    .Q(dsp_join_kb_26_TMR_1[6]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52657.11-52663.2" *)
  FD1P3IX \main_basesoc_tx_phase[6]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(N_17827_0_TMR_2),
    .Q(dsp_join_kb_26_TMR_2[6]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52664.11-52670.2" *)
  FD1P3IX \main_basesoc_tx_phase[7]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(N_17829_0_TMR_0),
    .Q(dsp_join_kb_26_TMR_0[7]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52664.11-52670.2" *)
  FD1P3IX \main_basesoc_tx_phase[7]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(N_17829_0_TMR_1),
    .Q(dsp_join_kb_26_TMR_1[7]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52664.11-52670.2" *)
  FD1P3IX \main_basesoc_tx_phase[7]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(N_17829_0_TMR_2),
    .Q(dsp_join_kb_26_TMR_2[7]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52671.11-52677.2" *)
  FD1P3IX \main_basesoc_tx_phase[8]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(N_17831_0_TMR_0),
    .Q(dsp_join_kb_26_TMR_0[8]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52671.11-52677.2" *)
  FD1P3IX \main_basesoc_tx_phase[8]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(N_17831_0_TMR_1),
    .Q(dsp_join_kb_26_TMR_1[8]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52671.11-52677.2" *)
  FD1P3IX \main_basesoc_tx_phase[8]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(N_17831_0_TMR_2),
    .Q(dsp_join_kb_26_TMR_2[8]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52678.11-52684.2" *)
  FD1P3IX \main_basesoc_tx_phase[9]_TMR_0  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_0),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_9_0_S0_TMR_0),
    .Q(dsp_join_kb_26_TMR_0[9]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52678.11-52684.2" *)
  FD1P3IX \main_basesoc_tx_phase[9]_TMR_1  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_1),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_9_0_S0_TMR_1),
    .Q(dsp_join_kb_26_TMR_1[9]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52678.11-52684.2" *)
  FD1P3IX \main_basesoc_tx_phase[9]_TMR_2  (
    .CD(builder_basesoc_rs232phytx_state_i_TMR_2),
    .CK(sys_clk),
    .D(un5_main_basesoc_tx_phase_cry_9_0_S0_TMR_2),
    .Q(dsp_join_kb_26_TMR_2[9]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51651.8-51657.2" *)
  LUT4 \main_basesoc_tx_phase_RNO[11]_TMR_0  (
    .A(builder_basesoc_rs232phytx_state_TMR_0),
    .B(un5_main_basesoc_tx_phase_cry_11_0_S0_TMR_0),
    .C(GND_0),
    .D(GND_0),
    .Z(N_17833_0_TMR_0)
  );
  defparam \main_basesoc_tx_phase_RNO[11]_TMR_0 .INIT = "0xDDDD";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51651.8-51657.2" *)
  LUT4 \main_basesoc_tx_phase_RNO[11]_TMR_1  (
    .A(builder_basesoc_rs232phytx_state_TMR_1),
    .B(un5_main_basesoc_tx_phase_cry_11_0_S0_TMR_1),
    .C(GND_0),
    .D(GND_0),
    .Z(N_17833_0_TMR_1)
  );
  defparam \main_basesoc_tx_phase_RNO[11]_TMR_1 .INIT = "0xDDDD";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51651.8-51657.2" *)
  LUT4 \main_basesoc_tx_phase_RNO[11]_TMR_2  (
    .A(builder_basesoc_rs232phytx_state_TMR_2),
    .B(un5_main_basesoc_tx_phase_cry_11_0_S0_TMR_2),
    .C(GND_0),
    .D(GND_0),
    .Z(N_17833_0_TMR_2)
  );
  defparam \main_basesoc_tx_phase_RNO[11]_TMR_2 .INIT = "0xDDDD";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51659.8-51665.2" *)
  LUT4 \main_basesoc_tx_phase_RNO[13]_TMR_0  (
    .A(builder_basesoc_rs232phytx_state_TMR_0),
    .B(un5_main_basesoc_tx_phase_cry_13_0_S0_TMR_0),
    .C(GND_0),
    .D(GND_0),
    .Z(N_17835_0_TMR_0)
  );
  defparam \main_basesoc_tx_phase_RNO[13]_TMR_0 .INIT = "0xDDDD";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51659.8-51665.2" *)
  LUT4 \main_basesoc_tx_phase_RNO[13]_TMR_1  (
    .A(builder_basesoc_rs232phytx_state_TMR_1),
    .B(un5_main_basesoc_tx_phase_cry_13_0_S0_TMR_1),
    .C(GND_0),
    .D(GND_0),
    .Z(N_17835_0_TMR_1)
  );
  defparam \main_basesoc_tx_phase_RNO[13]_TMR_1 .INIT = "0xDDDD";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51659.8-51665.2" *)
  LUT4 \main_basesoc_tx_phase_RNO[13]_TMR_2  (
    .A(builder_basesoc_rs232phytx_state_TMR_2),
    .B(un5_main_basesoc_tx_phase_cry_13_0_S0_TMR_2),
    .C(GND_0),
    .D(GND_0),
    .Z(N_17835_0_TMR_2)
  );
  defparam \main_basesoc_tx_phase_RNO[13]_TMR_2 .INIT = "0xDDDD";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51579.8-51585.2" *)
  LUT4 \main_basesoc_tx_phase_RNO[15]_TMR_0  (
    .A(builder_basesoc_rs232phytx_state_TMR_0),
    .B(un5_main_basesoc_tx_phase_cry_15_0_S0_TMR_0),
    .C(GND_0),
    .D(GND_0),
    .Z(N_17815_0_TMR_0)
  );
  defparam \main_basesoc_tx_phase_RNO[15]_TMR_0 .INIT = "0xDDDD";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51579.8-51585.2" *)
  LUT4 \main_basesoc_tx_phase_RNO[15]_TMR_1  (
    .A(builder_basesoc_rs232phytx_state_TMR_1),
    .B(un5_main_basesoc_tx_phase_cry_15_0_S0_TMR_1),
    .C(GND_0),
    .D(GND_0),
    .Z(N_17815_0_TMR_1)
  );
  defparam \main_basesoc_tx_phase_RNO[15]_TMR_1 .INIT = "0xDDDD";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51579.8-51585.2" *)
  LUT4 \main_basesoc_tx_phase_RNO[15]_TMR_2  (
    .A(builder_basesoc_rs232phytx_state_TMR_2),
    .B(un5_main_basesoc_tx_phase_cry_15_0_S0_TMR_2),
    .C(GND_0),
    .D(GND_0),
    .Z(N_17815_0_TMR_2)
  );
  defparam \main_basesoc_tx_phase_RNO[15]_TMR_2 .INIT = "0xDDDD";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51587.8-51593.2" *)
  LUT4 \main_basesoc_tx_phase_RNO[18]_TMR_0  (
    .A(builder_basesoc_rs232phytx_state_TMR_0),
    .B(un5_main_basesoc_tx_phase_cry_17_0_S1_TMR_0),
    .C(GND_0),
    .D(GND_0),
    .Z(N_17817_0_TMR_0)
  );
  defparam \main_basesoc_tx_phase_RNO[18]_TMR_0 .INIT = "0xDDDD";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51587.8-51593.2" *)
  LUT4 \main_basesoc_tx_phase_RNO[18]_TMR_1  (
    .A(builder_basesoc_rs232phytx_state_TMR_1),
    .B(un5_main_basesoc_tx_phase_cry_17_0_S1_TMR_1),
    .C(GND_0),
    .D(GND_0),
    .Z(N_17817_0_TMR_1)
  );
  defparam \main_basesoc_tx_phase_RNO[18]_TMR_1 .INIT = "0xDDDD";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51587.8-51593.2" *)
  LUT4 \main_basesoc_tx_phase_RNO[18]_TMR_2  (
    .A(builder_basesoc_rs232phytx_state_TMR_2),
    .B(un5_main_basesoc_tx_phase_cry_17_0_S1_TMR_2),
    .C(GND_0),
    .D(GND_0),
    .Z(N_17817_0_TMR_2)
  );
  defparam \main_basesoc_tx_phase_RNO[18]_TMR_2 .INIT = "0xDDDD";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51595.8-51601.2" *)
  LUT4 \main_basesoc_tx_phase_RNO[21]_TMR_0  (
    .A(builder_basesoc_rs232phytx_state_TMR_0),
    .B(un5_main_basesoc_tx_phase_cry_21_0_S0_TMR_0),
    .C(GND_0),
    .D(GND_0),
    .Z(N_17819_0_TMR_0)
  );
  defparam \main_basesoc_tx_phase_RNO[21]_TMR_0 .INIT = "0xDDDD";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51595.8-51601.2" *)
  LUT4 \main_basesoc_tx_phase_RNO[21]_TMR_1  (
    .A(builder_basesoc_rs232phytx_state_TMR_1),
    .B(un5_main_basesoc_tx_phase_cry_21_0_S0_TMR_1),
    .C(GND_0),
    .D(GND_0),
    .Z(N_17819_0_TMR_1)
  );
  defparam \main_basesoc_tx_phase_RNO[21]_TMR_1 .INIT = "0xDDDD";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51595.8-51601.2" *)
  LUT4 \main_basesoc_tx_phase_RNO[21]_TMR_2  (
    .A(builder_basesoc_rs232phytx_state_TMR_2),
    .B(un5_main_basesoc_tx_phase_cry_21_0_S0_TMR_2),
    .C(GND_0),
    .D(GND_0),
    .Z(N_17819_0_TMR_2)
  );
  defparam \main_basesoc_tx_phase_RNO[21]_TMR_2 .INIT = "0xDDDD";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51603.8-51609.2" *)
  LUT4 \main_basesoc_tx_phase_RNO[22]_TMR_0  (
    .A(builder_basesoc_rs232phytx_state_TMR_0),
    .B(un5_main_basesoc_tx_phase_cry_21_0_S1_TMR_0),
    .C(GND_0),
    .D(GND_0),
    .Z(N_17821_0_TMR_0)
  );
  defparam \main_basesoc_tx_phase_RNO[22]_TMR_0 .INIT = "0xDDDD";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51603.8-51609.2" *)
  LUT4 \main_basesoc_tx_phase_RNO[22]_TMR_1  (
    .A(builder_basesoc_rs232phytx_state_TMR_1),
    .B(un5_main_basesoc_tx_phase_cry_21_0_S1_TMR_1),
    .C(GND_0),
    .D(GND_0),
    .Z(N_17821_0_TMR_1)
  );
  defparam \main_basesoc_tx_phase_RNO[22]_TMR_1 .INIT = "0xDDDD";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51603.8-51609.2" *)
  LUT4 \main_basesoc_tx_phase_RNO[22]_TMR_2  (
    .A(builder_basesoc_rs232phytx_state_TMR_2),
    .B(un5_main_basesoc_tx_phase_cry_21_0_S1_TMR_2),
    .C(GND_0),
    .D(GND_0),
    .Z(N_17821_0_TMR_2)
  );
  defparam \main_basesoc_tx_phase_RNO[22]_TMR_2 .INIT = "0xDDDD";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51611.8-51617.2" *)
  LUT4 \main_basesoc_tx_phase_RNO[2]_TMR_0  (
    .A(builder_basesoc_rs232phytx_state_TMR_0),
    .B(un5_main_basesoc_tx_phase_cry_1_0_S1_TMR_0),
    .C(GND_0),
    .D(GND_0),
    .Z(N_17823_0_TMR_0)
  );
  defparam \main_basesoc_tx_phase_RNO[2]_TMR_0 .INIT = "0xDDDD";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51611.8-51617.2" *)
  LUT4 \main_basesoc_tx_phase_RNO[2]_TMR_1  (
    .A(builder_basesoc_rs232phytx_state_TMR_1),
    .B(un5_main_basesoc_tx_phase_cry_1_0_S1_TMR_1),
    .C(GND_0),
    .D(GND_0),
    .Z(N_17823_0_TMR_1)
  );
  defparam \main_basesoc_tx_phase_RNO[2]_TMR_1 .INIT = "0xDDDD";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51611.8-51617.2" *)
  LUT4 \main_basesoc_tx_phase_RNO[2]_TMR_2  (
    .A(builder_basesoc_rs232phytx_state_TMR_2),
    .B(un5_main_basesoc_tx_phase_cry_1_0_S1_TMR_2),
    .C(GND_0),
    .D(GND_0),
    .Z(N_17823_0_TMR_2)
  );
  defparam \main_basesoc_tx_phase_RNO[2]_TMR_2 .INIT = "0xDDDD";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51619.8-51625.2" *)
  LUT4 \main_basesoc_tx_phase_RNO[3]_TMR_0  (
    .A(builder_basesoc_rs232phytx_state_TMR_0),
    .B(un5_main_basesoc_tx_phase_cry_3_0_S0_TMR_0),
    .C(GND_0),
    .D(GND_0),
    .Z(N_17825_0_TMR_0)
  );
  defparam \main_basesoc_tx_phase_RNO[3]_TMR_0 .INIT = "0xDDDD";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51619.8-51625.2" *)
  LUT4 \main_basesoc_tx_phase_RNO[3]_TMR_1  (
    .A(builder_basesoc_rs232phytx_state_TMR_1),
    .B(un5_main_basesoc_tx_phase_cry_3_0_S0_TMR_1),
    .C(GND_0),
    .D(GND_0),
    .Z(N_17825_0_TMR_1)
  );
  defparam \main_basesoc_tx_phase_RNO[3]_TMR_1 .INIT = "0xDDDD";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51619.8-51625.2" *)
  LUT4 \main_basesoc_tx_phase_RNO[3]_TMR_2  (
    .A(builder_basesoc_rs232phytx_state_TMR_2),
    .B(un5_main_basesoc_tx_phase_cry_3_0_S0_TMR_2),
    .C(GND_0),
    .D(GND_0),
    .Z(N_17825_0_TMR_2)
  );
  defparam \main_basesoc_tx_phase_RNO[3]_TMR_2 .INIT = "0xDDDD";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51627.8-51633.2" *)
  LUT4 \main_basesoc_tx_phase_RNO[6]_TMR_0  (
    .A(builder_basesoc_rs232phytx_state_TMR_0),
    .B(un5_main_basesoc_tx_phase_cry_5_0_S1_TMR_0),
    .C(GND_0),
    .D(GND_0),
    .Z(N_17827_0_TMR_0)
  );
  defparam \main_basesoc_tx_phase_RNO[6]_TMR_0 .INIT = "0xDDDD";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51627.8-51633.2" *)
  LUT4 \main_basesoc_tx_phase_RNO[6]_TMR_1  (
    .A(builder_basesoc_rs232phytx_state_TMR_1),
    .B(un5_main_basesoc_tx_phase_cry_5_0_S1_TMR_1),
    .C(GND_0),
    .D(GND_0),
    .Z(N_17827_0_TMR_1)
  );
  defparam \main_basesoc_tx_phase_RNO[6]_TMR_1 .INIT = "0xDDDD";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51627.8-51633.2" *)
  LUT4 \main_basesoc_tx_phase_RNO[6]_TMR_2  (
    .A(builder_basesoc_rs232phytx_state_TMR_2),
    .B(un5_main_basesoc_tx_phase_cry_5_0_S1_TMR_2),
    .C(GND_0),
    .D(GND_0),
    .Z(N_17827_0_TMR_2)
  );
  defparam \main_basesoc_tx_phase_RNO[6]_TMR_2 .INIT = "0xDDDD";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51635.8-51641.2" *)
  LUT4 \main_basesoc_tx_phase_RNO[7]_TMR_0  (
    .A(builder_basesoc_rs232phytx_state_TMR_0),
    .B(un5_main_basesoc_tx_phase_cry_7_0_S0_TMR_0),
    .C(GND_0),
    .D(GND_0),
    .Z(N_17829_0_TMR_0)
  );
  defparam \main_basesoc_tx_phase_RNO[7]_TMR_0 .INIT = "0xDDDD";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51635.8-51641.2" *)
  LUT4 \main_basesoc_tx_phase_RNO[7]_TMR_1  (
    .A(builder_basesoc_rs232phytx_state_TMR_1),
    .B(un5_main_basesoc_tx_phase_cry_7_0_S0_TMR_1),
    .C(GND_0),
    .D(GND_0),
    .Z(N_17829_0_TMR_1)
  );
  defparam \main_basesoc_tx_phase_RNO[7]_TMR_1 .INIT = "0xDDDD";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51635.8-51641.2" *)
  LUT4 \main_basesoc_tx_phase_RNO[7]_TMR_2  (
    .A(builder_basesoc_rs232phytx_state_TMR_2),
    .B(un5_main_basesoc_tx_phase_cry_7_0_S0_TMR_2),
    .C(GND_0),
    .D(GND_0),
    .Z(N_17829_0_TMR_2)
  );
  defparam \main_basesoc_tx_phase_RNO[7]_TMR_2 .INIT = "0xDDDD";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51643.8-51649.2" *)
  LUT4 \main_basesoc_tx_phase_RNO[8]_TMR_0  (
    .A(builder_basesoc_rs232phytx_state_TMR_0),
    .B(un5_main_basesoc_tx_phase_cry_7_0_S1_TMR_0),
    .C(GND_0),
    .D(GND_0),
    .Z(N_17831_0_TMR_0)
  );
  defparam \main_basesoc_tx_phase_RNO[8]_TMR_0 .INIT = "0xDDDD";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51643.8-51649.2" *)
  LUT4 \main_basesoc_tx_phase_RNO[8]_TMR_1  (
    .A(builder_basesoc_rs232phytx_state_TMR_1),
    .B(un5_main_basesoc_tx_phase_cry_7_0_S1_TMR_1),
    .C(GND_0),
    .D(GND_0),
    .Z(N_17831_0_TMR_1)
  );
  defparam \main_basesoc_tx_phase_RNO[8]_TMR_1 .INIT = "0xDDDD";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51643.8-51649.2" *)
  LUT4 \main_basesoc_tx_phase_RNO[8]_TMR_2  (
    .A(builder_basesoc_rs232phytx_state_TMR_2),
    .B(un5_main_basesoc_tx_phase_cry_7_0_S1_TMR_2),
    .C(GND_0),
    .D(GND_0),
    .Z(N_17831_0_TMR_2)
  );
  defparam \main_basesoc_tx_phase_RNO[8]_TMR_2 .INIT = "0xDDDD";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52615.11-52621.2" *)
  FD1P3IX \main_basesoc_tx_phase_mod[0]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_tx_phase_mod_RNO_TMR_0),
    .Q(dsp_join_kb_26_TMR_0[0]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52615.11-52621.2" *)
  FD1P3IX \main_basesoc_tx_phase_mod[0]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_tx_phase_mod_RNO_TMR_1),
    .Q(dsp_join_kb_26_TMR_1[0]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52615.11-52621.2" *)
  FD1P3IX \main_basesoc_tx_phase_mod[0]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_tx_phase_mod_RNO_TMR_2),
    .Q(dsp_join_kb_26_TMR_2[0]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56210.8-56216.2" *)
  LUT4 \main_basesoc_tx_phase_mod_RNO_cZ[0]_TMR_0  (
    .A(builder_basesoc_rs232phytx_state_TMR_0),
    .B(dsp_join_kb_26_TMR_0[0]),
    .C(GND_0),
    .D(GND_0),
    .Z(main_basesoc_tx_phase_mod_RNO_TMR_0)
  );
  defparam \main_basesoc_tx_phase_mod_RNO_cZ[0]_TMR_0 .INIT = "0x7777";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56210.8-56216.2" *)
  LUT4 \main_basesoc_tx_phase_mod_RNO_cZ[0]_TMR_1  (
    .A(builder_basesoc_rs232phytx_state_TMR_1),
    .B(dsp_join_kb_26_TMR_1[0]),
    .C(GND_0),
    .D(GND_0),
    .Z(main_basesoc_tx_phase_mod_RNO_TMR_1)
  );
  defparam \main_basesoc_tx_phase_mod_RNO_cZ[0]_TMR_1 .INIT = "0x7777";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56210.8-56216.2" *)
  LUT4 \main_basesoc_tx_phase_mod_RNO_cZ[0]_TMR_2  (
    .A(builder_basesoc_rs232phytx_state_TMR_2),
    .B(dsp_join_kb_26_TMR_2[0]),
    .C(GND_0),
    .D(GND_0),
    .Z(main_basesoc_tx_phase_mod_RNO_TMR_2)
  );
  defparam \main_basesoc_tx_phase_mod_RNO_cZ[0]_TMR_2 .INIT = "0x7777";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52608.11-52614.2" *)
  FD1P3IX main_basesoc_tx_tick_reg_TMR_0 (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(main_basesoc_tx_tick_0_TMR_0),
    .Q(main_basesoc_tx_tick_TMR_0),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52608.11-52614.2" *)
  FD1P3IX main_basesoc_tx_tick_reg_TMR_1 (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(main_basesoc_tx_tick_0_TMR_1),
    .Q(main_basesoc_tx_tick_TMR_1),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52608.11-52614.2" *)
  FD1P3IX main_basesoc_tx_tick_reg_TMR_2 (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(main_basesoc_tx_tick_0_TMR_2),
    .Q(main_basesoc_tx_tick_TMR_2),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52594.11-52600.2" *)
  FD1P3IX \main_basesoc_uart_enable_storage_reg[0]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[0]),
    .Q(main_basesoc_uart_enable_storage_TMR_0[0]),
    .SP(builder_csr_bankarray_csrbank3_ev_enable0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52594.11-52600.2" *)
  FD1P3IX \main_basesoc_uart_enable_storage_reg[0]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[0]),
    .Q(main_basesoc_uart_enable_storage_TMR_1[0]),
    .SP(builder_csr_bankarray_csrbank3_ev_enable0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52594.11-52600.2" *)
  FD1P3IX \main_basesoc_uart_enable_storage_reg[0]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[0]),
    .Q(main_basesoc_uart_enable_storage_TMR_2[0]),
    .SP(builder_csr_bankarray_csrbank3_ev_enable0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52601.11-52607.2" *)
  FD1P3IX \main_basesoc_uart_enable_storage_reg[1]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[1]),
    .Q(main_basesoc_uart_enable_storage_TMR_0[1]),
    .SP(builder_csr_bankarray_csrbank3_ev_enable0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52601.11-52607.2" *)
  FD1P3IX \main_basesoc_uart_enable_storage_reg[1]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[1]),
    .Q(main_basesoc_uart_enable_storage_TMR_1[1]),
    .SP(builder_csr_bankarray_csrbank3_ev_enable0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52601.11-52607.2" *)
  FD1P3IX \main_basesoc_uart_enable_storage_reg[1]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[1]),
    .Q(main_basesoc_uart_enable_storage_TMR_2[1]),
    .SP(builder_csr_bankarray_csrbank3_ev_enable0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52580.11-52586.2" *)
  FD1P3IX \main_basesoc_uart_pending_r_reg[0]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[0]),
    .Q(main_basesoc_uart_pending_r_TMR_0[0]),
    .SP(builder_csr_bankarray_csrbank3_ev_pending_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52580.11-52586.2" *)
  FD1P3IX \main_basesoc_uart_pending_r_reg[0]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[0]),
    .Q(main_basesoc_uart_pending_r_TMR_1[0]),
    .SP(builder_csr_bankarray_csrbank3_ev_pending_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52580.11-52586.2" *)
  FD1P3IX \main_basesoc_uart_pending_r_reg[0]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[0]),
    .Q(main_basesoc_uart_pending_r_TMR_2[0]),
    .SP(builder_csr_bankarray_csrbank3_ev_pending_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52587.11-52593.2" *)
  FD1P3IX \main_basesoc_uart_pending_r_reg[1]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[1]),
    .Q(main_basesoc_uart_pending_r_TMR_0[1]),
    .SP(builder_csr_bankarray_csrbank3_ev_pending_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52587.11-52593.2" *)
  FD1P3IX \main_basesoc_uart_pending_r_reg[1]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[1]),
    .Q(main_basesoc_uart_pending_r_TMR_1[1]),
    .SP(builder_csr_bankarray_csrbank3_ev_pending_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52587.11-52593.2" *)
  FD1P3IX \main_basesoc_uart_pending_r_reg[1]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[1]),
    .Q(main_basesoc_uart_pending_r_TMR_2[1]),
    .SP(builder_csr_bankarray_csrbank3_ev_pending_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52573.11-52579.2" *)
  FD1P3IX main_basesoc_uart_pending_re_reg_TMR_0 (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_uart_pending_r_0_sqmuxa_TMR_0),
    .Q(main_basesoc_uart_pending_re_TMR_0),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52573.11-52579.2" *)
  FD1P3IX main_basesoc_uart_pending_re_reg_TMR_1 (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_uart_pending_r_0_sqmuxa_TMR_1),
    .Q(main_basesoc_uart_pending_re_TMR_1),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52573.11-52579.2" *)
  FD1P3IX main_basesoc_uart_pending_re_reg_TMR_2 (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_uart_pending_r_0_sqmuxa_TMR_2),
    .Q(main_basesoc_uart_pending_re_TMR_2),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51362.8-51368.2" *)
  LUT4 \main_basesoc_uart_rx_fifo_consume_RNO_cZ[2]_TMR_0  (
    .A(main_basesoc_uart_rx_fifo_consume_TMR_0[2]),
    .B(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_0),
    .C(main_basesoc_uart_rx_fifo_consume_TMR_0[1]),
    .D(main_basesoc_uart_rx_fifo_consume_TMR_0[0]),
    .Z(main_basesoc_uart_rx_fifo_consume_RNO_TMR_0)
  );
  defparam \main_basesoc_uart_rx_fifo_consume_RNO_cZ[2]_TMR_0 .INIT = "0x6AAA";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51362.8-51368.2" *)
  LUT4 \main_basesoc_uart_rx_fifo_consume_RNO_cZ[2]_TMR_1  (
    .A(main_basesoc_uart_rx_fifo_consume_TMR_1[2]),
    .B(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_1),
    .C(main_basesoc_uart_rx_fifo_consume_TMR_1[1]),
    .D(main_basesoc_uart_rx_fifo_consume_TMR_1[0]),
    .Z(main_basesoc_uart_rx_fifo_consume_RNO_TMR_1)
  );
  defparam \main_basesoc_uart_rx_fifo_consume_RNO_cZ[2]_TMR_1 .INIT = "0x6AAA";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51362.8-51368.2" *)
  LUT4 \main_basesoc_uart_rx_fifo_consume_RNO_cZ[2]_TMR_2  (
    .A(main_basesoc_uart_rx_fifo_consume_TMR_2[2]),
    .B(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_2),
    .C(main_basesoc_uart_rx_fifo_consume_TMR_2[1]),
    .D(main_basesoc_uart_rx_fifo_consume_TMR_2[0]),
    .Z(main_basesoc_uart_rx_fifo_consume_RNO_TMR_2)
  );
  defparam \main_basesoc_uart_rx_fifo_consume_RNO_cZ[2]_TMR_2 .INIT = "0x6AAA";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52545.11-52551.2" *)
  FD1P3IX \main_basesoc_uart_rx_fifo_consume_reg[0]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_rx_fifo_consume_axbxc0_TMR_0),
    .Q(main_basesoc_uart_rx_fifo_consume_TMR_0[0]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52545.11-52551.2" *)
  FD1P3IX \main_basesoc_uart_rx_fifo_consume_reg[0]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_rx_fifo_consume_axbxc0_TMR_1),
    .Q(main_basesoc_uart_rx_fifo_consume_TMR_1[0]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52545.11-52551.2" *)
  FD1P3IX \main_basesoc_uart_rx_fifo_consume_reg[0]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_rx_fifo_consume_axbxc0_TMR_2),
    .Q(main_basesoc_uart_rx_fifo_consume_TMR_2[0]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52552.11-52558.2" *)
  FD1P3IX \main_basesoc_uart_rx_fifo_consume_reg[1]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_rx_fifo_consume_axbxc1_TMR_0),
    .Q(main_basesoc_uart_rx_fifo_consume_TMR_0[1]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52552.11-52558.2" *)
  FD1P3IX \main_basesoc_uart_rx_fifo_consume_reg[1]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_rx_fifo_consume_axbxc1_TMR_1),
    .Q(main_basesoc_uart_rx_fifo_consume_TMR_1[1]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52552.11-52558.2" *)
  FD1P3IX \main_basesoc_uart_rx_fifo_consume_reg[1]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_rx_fifo_consume_axbxc1_TMR_2),
    .Q(main_basesoc_uart_rx_fifo_consume_TMR_2[1]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52559.11-52565.2" *)
  FD1P3IX \main_basesoc_uart_rx_fifo_consume_reg[2]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(main_basesoc_uart_rx_fifo_consume_RNO_TMR_0),
    .Q(main_basesoc_uart_rx_fifo_consume_TMR_0[2]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52559.11-52565.2" *)
  FD1P3IX \main_basesoc_uart_rx_fifo_consume_reg[2]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(main_basesoc_uart_rx_fifo_consume_RNO_TMR_1),
    .Q(main_basesoc_uart_rx_fifo_consume_TMR_1[2]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52559.11-52565.2" *)
  FD1P3IX \main_basesoc_uart_rx_fifo_consume_reg[2]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(main_basesoc_uart_rx_fifo_consume_RNO_TMR_2),
    .Q(main_basesoc_uart_rx_fifo_consume_TMR_2[2]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52566.11-52572.2" *)
  FD1P3IX \main_basesoc_uart_rx_fifo_consume_reg[3]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_rx_fifo_consume_axbxc3_TMR_0),
    .Q(main_basesoc_uart_rx_fifo_consume_TMR_0[3]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52566.11-52572.2" *)
  FD1P3IX \main_basesoc_uart_rx_fifo_consume_reg[3]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_rx_fifo_consume_axbxc3_TMR_1),
    .Q(main_basesoc_uart_rx_fifo_consume_TMR_1[3]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52566.11-52572.2" *)
  FD1P3IX \main_basesoc_uart_rx_fifo_consume_reg[3]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_rx_fifo_consume_axbxc3_TMR_2),
    .Q(main_basesoc_uart_rx_fifo_consume_TMR_2[3]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52524.11-52530.2" *)
  FD1P3IX \main_basesoc_uart_rx_fifo_level0_0_mod[0]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_uart_rx_fifo_level0_0_mod_RNO_TMR_0),
    .Q(un1_main_basesoc_uart_rx_fifo_level0_scalar_TMR_0),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52524.11-52530.2" *)
  FD1P3IX \main_basesoc_uart_rx_fifo_level0_0_mod[0]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_uart_rx_fifo_level0_0_mod_RNO_TMR_1),
    .Q(un1_main_basesoc_uart_rx_fifo_level0_scalar_TMR_1),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52524.11-52530.2" *)
  FD1P3IX \main_basesoc_uart_rx_fifo_level0_0_mod[0]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_uart_rx_fifo_level0_0_mod_RNO_TMR_2),
    .Q(un1_main_basesoc_uart_rx_fifo_level0_scalar_TMR_2),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52531.11-52537.2" *)
  FD1P3IX \main_basesoc_uart_rx_fifo_level0_0_mod[2]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_rx_fifo_level0_TMR_0[2]),
    .Q(un1_main_basesoc_uart_rx_fifo_level0_0_TMR_0[2]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52531.11-52537.2" *)
  FD1P3IX \main_basesoc_uart_rx_fifo_level0_0_mod[2]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_rx_fifo_level0_TMR_1[2]),
    .Q(un1_main_basesoc_uart_rx_fifo_level0_0_TMR_1[2]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52531.11-52537.2" *)
  FD1P3IX \main_basesoc_uart_rx_fifo_level0_0_mod[2]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_rx_fifo_level0_TMR_2[2]),
    .Q(un1_main_basesoc_uart_rx_fifo_level0_0_TMR_2[2]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52538.11-52544.2" *)
  FD1P3IX \main_basesoc_uart_rx_fifo_level0_0_mod[4]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_rx_fifo_level0_TMR_0[4]),
    .Q(un1_main_basesoc_uart_rx_fifo_level0_0_TMR_0[4]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52538.11-52544.2" *)
  FD1P3IX \main_basesoc_uart_rx_fifo_level0_0_mod[4]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_rx_fifo_level0_TMR_1[4]),
    .Q(un1_main_basesoc_uart_rx_fifo_level0_0_TMR_1[4]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52538.11-52544.2" *)
  FD1P3IX \main_basesoc_uart_rx_fifo_level0_0_mod[4]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_rx_fifo_level0_TMR_2[4]),
    .Q(un1_main_basesoc_uart_rx_fifo_level0_0_TMR_2[4]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55629.8-55635.2" *)
  LUT4 \main_basesoc_uart_rx_fifo_level0_0_mod_RNO_cZ[0]_TMR_0  (
    .A(sys_rst_TMR_0),
    .B(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_0),
    .C(main_basesoc_uart_rx_fifo_wrport_we_TMR_0),
    .D(un1_main_basesoc_uart_rx_fifo_level0_scalar_TMR_0),
    .Z(main_basesoc_uart_rx_fifo_level0_0_mod_RNO_TMR_0)
  );
  defparam \main_basesoc_uart_rx_fifo_level0_0_mod_RNO_cZ[0]_TMR_0 .INIT = "0x4114";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55629.8-55635.2" *)
  LUT4 \main_basesoc_uart_rx_fifo_level0_0_mod_RNO_cZ[0]_TMR_1  (
    .A(sys_rst_TMR_1),
    .B(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_1),
    .C(main_basesoc_uart_rx_fifo_wrport_we_TMR_1),
    .D(un1_main_basesoc_uart_rx_fifo_level0_scalar_TMR_1),
    .Z(main_basesoc_uart_rx_fifo_level0_0_mod_RNO_TMR_1)
  );
  defparam \main_basesoc_uart_rx_fifo_level0_0_mod_RNO_cZ[0]_TMR_1 .INIT = "0x4114";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55629.8-55635.2" *)
  LUT4 \main_basesoc_uart_rx_fifo_level0_0_mod_RNO_cZ[0]_TMR_2  (
    .A(sys_rst_TMR_2),
    .B(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_2),
    .C(main_basesoc_uart_rx_fifo_wrport_we_TMR_2),
    .D(un1_main_basesoc_uart_rx_fifo_level0_scalar_TMR_2),
    .Z(main_basesoc_uart_rx_fifo_level0_0_mod_RNO_TMR_2)
  );
  defparam \main_basesoc_uart_rx_fifo_level0_0_mod_RNO_cZ[0]_TMR_2 .INIT = "0x4114";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52510.11-52516.2" *)
  FD1P3IX \main_basesoc_uart_rx_fifo_level0_mod[1]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_rx_fifo_level0_TMR_0[1]),
    .Q(un1_main_basesoc_uart_rx_fifo_level0_0_TMR_0[1]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52510.11-52516.2" *)
  FD1P3IX \main_basesoc_uart_rx_fifo_level0_mod[1]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_rx_fifo_level0_TMR_1[1]),
    .Q(un1_main_basesoc_uart_rx_fifo_level0_0_TMR_1[1]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52510.11-52516.2" *)
  FD1P3IX \main_basesoc_uart_rx_fifo_level0_mod[1]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_rx_fifo_level0_TMR_2[1]),
    .Q(un1_main_basesoc_uart_rx_fifo_level0_0_TMR_2[1]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52517.11-52523.2" *)
  FD1P3IX \main_basesoc_uart_rx_fifo_level0_mod[3]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_rx_fifo_level0_TMR_0[3]),
    .Q(un1_main_basesoc_uart_rx_fifo_level0_0_TMR_0[3]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52517.11-52523.2" *)
  FD1P3IX \main_basesoc_uart_rx_fifo_level0_mod[3]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_rx_fifo_level0_TMR_1[3]),
    .Q(un1_main_basesoc_uart_rx_fifo_level0_0_TMR_1[3]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52517.11-52523.2" *)
  FD1P3IX \main_basesoc_uart_rx_fifo_level0_mod[3]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_rx_fifo_level0_TMR_2[3]),
    .Q(un1_main_basesoc_uart_rx_fifo_level0_0_TMR_2[3]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51371.8-51377.2" *)
  LUT4 \main_basesoc_uart_rx_fifo_produce_RNO_cZ[2]_TMR_0  (
    .A(main_basesoc_uart_rx_fifo_produce_TMR_0[2]),
    .B(main_basesoc_uart_rx_fifo_wrport_we_TMR_0),
    .C(main_basesoc_uart_rx_fifo_produce_TMR_0[1]),
    .D(main_basesoc_uart_rx_fifo_produce_TMR_0[0]),
    .Z(main_basesoc_uart_rx_fifo_produce_RNO_TMR_0)
  );
  defparam \main_basesoc_uart_rx_fifo_produce_RNO_cZ[2]_TMR_0 .INIT = "0x6AAA";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51371.8-51377.2" *)
  LUT4 \main_basesoc_uart_rx_fifo_produce_RNO_cZ[2]_TMR_1  (
    .A(main_basesoc_uart_rx_fifo_produce_TMR_1[2]),
    .B(main_basesoc_uart_rx_fifo_wrport_we_TMR_1),
    .C(main_basesoc_uart_rx_fifo_produce_TMR_1[1]),
    .D(main_basesoc_uart_rx_fifo_produce_TMR_1[0]),
    .Z(main_basesoc_uart_rx_fifo_produce_RNO_TMR_1)
  );
  defparam \main_basesoc_uart_rx_fifo_produce_RNO_cZ[2]_TMR_1 .INIT = "0x6AAA";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51371.8-51377.2" *)
  LUT4 \main_basesoc_uart_rx_fifo_produce_RNO_cZ[2]_TMR_2  (
    .A(main_basesoc_uart_rx_fifo_produce_TMR_2[2]),
    .B(main_basesoc_uart_rx_fifo_wrport_we_TMR_2),
    .C(main_basesoc_uart_rx_fifo_produce_TMR_2[1]),
    .D(main_basesoc_uart_rx_fifo_produce_TMR_2[0]),
    .Z(main_basesoc_uart_rx_fifo_produce_RNO_TMR_2)
  );
  defparam \main_basesoc_uart_rx_fifo_produce_RNO_cZ[2]_TMR_2 .INIT = "0x6AAA";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52482.11-52488.2" *)
  FD1P3IX \main_basesoc_uart_rx_fifo_produce_reg[0]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_rx_fifo_produce_axbxc0_TMR_0),
    .Q(main_basesoc_uart_rx_fifo_produce_TMR_0[0]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52482.11-52488.2" *)
  FD1P3IX \main_basesoc_uart_rx_fifo_produce_reg[0]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_rx_fifo_produce_axbxc0_TMR_1),
    .Q(main_basesoc_uart_rx_fifo_produce_TMR_1[0]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52482.11-52488.2" *)
  FD1P3IX \main_basesoc_uart_rx_fifo_produce_reg[0]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_rx_fifo_produce_axbxc0_TMR_2),
    .Q(main_basesoc_uart_rx_fifo_produce_TMR_2[0]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52489.11-52495.2" *)
  FD1P3IX \main_basesoc_uart_rx_fifo_produce_reg[1]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_rx_fifo_produce_axbxc1_TMR_0),
    .Q(main_basesoc_uart_rx_fifo_produce_TMR_0[1]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52489.11-52495.2" *)
  FD1P3IX \main_basesoc_uart_rx_fifo_produce_reg[1]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_rx_fifo_produce_axbxc1_TMR_1),
    .Q(main_basesoc_uart_rx_fifo_produce_TMR_1[1]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52489.11-52495.2" *)
  FD1P3IX \main_basesoc_uart_rx_fifo_produce_reg[1]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_rx_fifo_produce_axbxc1_TMR_2),
    .Q(main_basesoc_uart_rx_fifo_produce_TMR_2[1]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52496.11-52502.2" *)
  FD1P3IX \main_basesoc_uart_rx_fifo_produce_reg[2]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(main_basesoc_uart_rx_fifo_produce_RNO_TMR_0),
    .Q(main_basesoc_uart_rx_fifo_produce_TMR_0[2]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52496.11-52502.2" *)
  FD1P3IX \main_basesoc_uart_rx_fifo_produce_reg[2]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(main_basesoc_uart_rx_fifo_produce_RNO_TMR_1),
    .Q(main_basesoc_uart_rx_fifo_produce_TMR_1[2]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52496.11-52502.2" *)
  FD1P3IX \main_basesoc_uart_rx_fifo_produce_reg[2]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(main_basesoc_uart_rx_fifo_produce_RNO_TMR_2),
    .Q(main_basesoc_uart_rx_fifo_produce_TMR_2[2]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52503.11-52509.2" *)
  FD1P3IX \main_basesoc_uart_rx_fifo_produce_reg[3]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_rx_fifo_produce_axbxc3_TMR_0),
    .Q(main_basesoc_uart_rx_fifo_produce_TMR_0[3]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52503.11-52509.2" *)
  FD1P3IX \main_basesoc_uart_rx_fifo_produce_reg[3]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_rx_fifo_produce_axbxc3_TMR_1),
    .Q(main_basesoc_uart_rx_fifo_produce_TMR_1[3]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52503.11-52509.2" *)
  FD1P3IX \main_basesoc_uart_rx_fifo_produce_reg[3]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_rx_fifo_produce_axbxc3_TMR_2),
    .Q(main_basesoc_uart_rx_fifo_produce_TMR_2[3]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52475.11-52481.2" *)
  FD1P3IX main_basesoc_uart_rx_fifo_readable_reg_TMR_0 (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(N_92_TMR_0),
    .Q(main_basesoc_uart_rx_fifo_readable_TMR_0),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52475.11-52481.2" *)
  FD1P3IX main_basesoc_uart_rx_fifo_readable_reg_TMR_1 (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(N_92_TMR_1),
    .Q(main_basesoc_uart_rx_fifo_readable_TMR_1),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52475.11-52481.2" *)
  FD1P3IX main_basesoc_uart_rx_fifo_readable_reg_TMR_2 (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(N_92_TMR_2),
    .Q(main_basesoc_uart_rx_fifo_readable_TMR_2),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52468.11-52474.2" *)
  FD1P3IX main_basesoc_uart_rx_pending_reg_TMR_0 (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(N_20_TMR_0),
    .Q(main_basesoc_uart_rx_pending_TMR_0),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52468.11-52474.2" *)
  FD1P3IX main_basesoc_uart_rx_pending_reg_TMR_1 (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(N_20_TMR_1),
    .Q(main_basesoc_uart_rx_pending_TMR_1),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52468.11-52474.2" *)
  FD1P3IX main_basesoc_uart_rx_pending_reg_TMR_2 (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(N_20_TMR_2),
    .Q(main_basesoc_uart_rx_pending_TMR_2),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52461.11-52467.2" *)
  FD1P3IX main_basesoc_uart_rx_trigger_d_reg_TMR_0 (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(main_basesoc_uart_rx_fifo_readable_TMR_0),
    .Q(main_basesoc_uart_rx_trigger_d_TMR_0),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52461.11-52467.2" *)
  FD1P3IX main_basesoc_uart_rx_trigger_d_reg_TMR_1 (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(main_basesoc_uart_rx_fifo_readable_TMR_1),
    .Q(main_basesoc_uart_rx_trigger_d_TMR_1),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52461.11-52467.2" *)
  FD1P3IX main_basesoc_uart_rx_trigger_d_reg_TMR_2 (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(main_basesoc_uart_rx_fifo_readable_TMR_2),
    .Q(main_basesoc_uart_rx_trigger_d_TMR_2),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51380.8-51386.2" *)
  LUT4 \main_basesoc_uart_tx_fifo_consume_RNO_cZ[2]_TMR_0  (
    .A(main_basesoc_uart_tx_fifo_consume_TMR_0[2]),
    .B(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_0),
    .C(main_basesoc_uart_tx_fifo_consume_TMR_0[1]),
    .D(main_basesoc_uart_tx_fifo_consume_TMR_0[0]),
    .Z(main_basesoc_uart_tx_fifo_consume_RNO_TMR_0)
  );
  defparam \main_basesoc_uart_tx_fifo_consume_RNO_cZ[2]_TMR_0 .INIT = "0x6AAA";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51380.8-51386.2" *)
  LUT4 \main_basesoc_uart_tx_fifo_consume_RNO_cZ[2]_TMR_1  (
    .A(main_basesoc_uart_tx_fifo_consume_TMR_1[2]),
    .B(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_1),
    .C(main_basesoc_uart_tx_fifo_consume_TMR_1[1]),
    .D(main_basesoc_uart_tx_fifo_consume_TMR_1[0]),
    .Z(main_basesoc_uart_tx_fifo_consume_RNO_TMR_1)
  );
  defparam \main_basesoc_uart_tx_fifo_consume_RNO_cZ[2]_TMR_1 .INIT = "0x6AAA";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51380.8-51386.2" *)
  LUT4 \main_basesoc_uart_tx_fifo_consume_RNO_cZ[2]_TMR_2  (
    .A(main_basesoc_uart_tx_fifo_consume_TMR_2[2]),
    .B(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_2),
    .C(main_basesoc_uart_tx_fifo_consume_TMR_2[1]),
    .D(main_basesoc_uart_tx_fifo_consume_TMR_2[0]),
    .Z(main_basesoc_uart_tx_fifo_consume_RNO_TMR_2)
  );
  defparam \main_basesoc_uart_tx_fifo_consume_RNO_cZ[2]_TMR_2 .INIT = "0x6AAA";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52433.11-52439.2" *)
  FD1P3IX \main_basesoc_uart_tx_fifo_consume_reg[0]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_tx_fifo_consume_axbxc0_TMR_0),
    .Q(main_basesoc_uart_tx_fifo_consume_TMR_0[0]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52433.11-52439.2" *)
  FD1P3IX \main_basesoc_uart_tx_fifo_consume_reg[0]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_tx_fifo_consume_axbxc0_TMR_1),
    .Q(main_basesoc_uart_tx_fifo_consume_TMR_1[0]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52433.11-52439.2" *)
  FD1P3IX \main_basesoc_uart_tx_fifo_consume_reg[0]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_tx_fifo_consume_axbxc0_TMR_2),
    .Q(main_basesoc_uart_tx_fifo_consume_TMR_2[0]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52440.11-52446.2" *)
  FD1P3IX \main_basesoc_uart_tx_fifo_consume_reg[1]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_tx_fifo_consume_axbxc1_TMR_0),
    .Q(main_basesoc_uart_tx_fifo_consume_TMR_0[1]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52440.11-52446.2" *)
  FD1P3IX \main_basesoc_uart_tx_fifo_consume_reg[1]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_tx_fifo_consume_axbxc1_TMR_1),
    .Q(main_basesoc_uart_tx_fifo_consume_TMR_1[1]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52440.11-52446.2" *)
  FD1P3IX \main_basesoc_uart_tx_fifo_consume_reg[1]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_tx_fifo_consume_axbxc1_TMR_2),
    .Q(main_basesoc_uart_tx_fifo_consume_TMR_2[1]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52447.11-52453.2" *)
  FD1P3IX \main_basesoc_uart_tx_fifo_consume_reg[2]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(main_basesoc_uart_tx_fifo_consume_RNO_TMR_0),
    .Q(main_basesoc_uart_tx_fifo_consume_TMR_0[2]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52447.11-52453.2" *)
  FD1P3IX \main_basesoc_uart_tx_fifo_consume_reg[2]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(main_basesoc_uart_tx_fifo_consume_RNO_TMR_1),
    .Q(main_basesoc_uart_tx_fifo_consume_TMR_1[2]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52447.11-52453.2" *)
  FD1P3IX \main_basesoc_uart_tx_fifo_consume_reg[2]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(main_basesoc_uart_tx_fifo_consume_RNO_TMR_2),
    .Q(main_basesoc_uart_tx_fifo_consume_TMR_2[2]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52454.11-52460.2" *)
  FD1P3IX \main_basesoc_uart_tx_fifo_consume_reg[3]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_tx_fifo_consume_axbxc3_TMR_0),
    .Q(main_basesoc_uart_tx_fifo_consume_TMR_0[3]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52454.11-52460.2" *)
  FD1P3IX \main_basesoc_uart_tx_fifo_consume_reg[3]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_tx_fifo_consume_axbxc3_TMR_1),
    .Q(main_basesoc_uart_tx_fifo_consume_TMR_1[3]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52454.11-52460.2" *)
  FD1P3IX \main_basesoc_uart_tx_fifo_consume_reg[3]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_tx_fifo_consume_axbxc3_TMR_2),
    .Q(main_basesoc_uart_tx_fifo_consume_TMR_2[3]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52412.11-52418.2" *)
  FD1P3IX \main_basesoc_uart_tx_fifo_level0_0_mod[0]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_uart_tx_fifo_level0_0_mod_RNO_TMR_0),
    .Q(un1_main_basesoc_uart_tx_fifo_level0_scalar_TMR_0),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52412.11-52418.2" *)
  FD1P3IX \main_basesoc_uart_tx_fifo_level0_0_mod[0]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_uart_tx_fifo_level0_0_mod_RNO_TMR_1),
    .Q(un1_main_basesoc_uart_tx_fifo_level0_scalar_TMR_1),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52412.11-52418.2" *)
  FD1P3IX \main_basesoc_uart_tx_fifo_level0_0_mod[0]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_basesoc_uart_tx_fifo_level0_0_mod_RNO_TMR_2),
    .Q(un1_main_basesoc_uart_tx_fifo_level0_scalar_TMR_2),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52419.11-52425.2" *)
  FD1P3IX \main_basesoc_uart_tx_fifo_level0_0_mod[2]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_tx_fifo_level0_TMR_0[2]),
    .Q(un1_main_basesoc_uart_tx_fifo_level0_0_TMR_0[2]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52419.11-52425.2" *)
  FD1P3IX \main_basesoc_uart_tx_fifo_level0_0_mod[2]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_tx_fifo_level0_TMR_1[2]),
    .Q(un1_main_basesoc_uart_tx_fifo_level0_0_TMR_1[2]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52419.11-52425.2" *)
  FD1P3IX \main_basesoc_uart_tx_fifo_level0_0_mod[2]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_tx_fifo_level0_TMR_2[2]),
    .Q(un1_main_basesoc_uart_tx_fifo_level0_0_TMR_2[2]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52426.11-52432.2" *)
  FD1P3IX \main_basesoc_uart_tx_fifo_level0_0_mod[4]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_tx_fifo_level0_TMR_0[4]),
    .Q(un1_main_basesoc_uart_tx_fifo_level0_0_TMR_0[4]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52426.11-52432.2" *)
  FD1P3IX \main_basesoc_uart_tx_fifo_level0_0_mod[4]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_tx_fifo_level0_TMR_1[4]),
    .Q(un1_main_basesoc_uart_tx_fifo_level0_0_TMR_1[4]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52426.11-52432.2" *)
  FD1P3IX \main_basesoc_uart_tx_fifo_level0_0_mod[4]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_tx_fifo_level0_TMR_2[4]),
    .Q(un1_main_basesoc_uart_tx_fifo_level0_0_TMR_2[4]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56335.8-56341.2" *)
  LUT4 \main_basesoc_uart_tx_fifo_level0_0_mod_RNIG0F3_cZ[0]_TMR_0  (
    .A(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_0),
    .B(un1_main_basesoc_uart_tx_fifo_level0_scalar_TMR_0),
    .C(GND_0),
    .D(GND_0),
    .Z(main_basesoc_uart_tx_fifo_level0_0_mod_RNIG0F3_TMR_0)
  );
  defparam \main_basesoc_uart_tx_fifo_level0_0_mod_RNIG0F3_cZ[0]_TMR_0 .INIT = "0x6666";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56335.8-56341.2" *)
  LUT4 \main_basesoc_uart_tx_fifo_level0_0_mod_RNIG0F3_cZ[0]_TMR_1  (
    .A(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_1),
    .B(un1_main_basesoc_uart_tx_fifo_level0_scalar_TMR_1),
    .C(GND_0),
    .D(GND_0),
    .Z(main_basesoc_uart_tx_fifo_level0_0_mod_RNIG0F3_TMR_1)
  );
  defparam \main_basesoc_uart_tx_fifo_level0_0_mod_RNIG0F3_cZ[0]_TMR_1 .INIT = "0x6666";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56335.8-56341.2" *)
  LUT4 \main_basesoc_uart_tx_fifo_level0_0_mod_RNIG0F3_cZ[0]_TMR_2  (
    .A(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_2),
    .B(un1_main_basesoc_uart_tx_fifo_level0_scalar_TMR_2),
    .C(GND_0),
    .D(GND_0),
    .Z(main_basesoc_uart_tx_fifo_level0_0_mod_RNIG0F3_TMR_2)
  );
  defparam \main_basesoc_uart_tx_fifo_level0_0_mod_RNIG0F3_cZ[0]_TMR_2 .INIT = "0x6666";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55586.8-55592.2" *)
  LUT4 \main_basesoc_uart_tx_fifo_level0_0_mod_RNO_cZ[0]_TMR_0  (
    .A(sys_rst_TMR_0),
    .B(un1_main_basesoc_uart_tx_fifo_level0_TMR_0[0]),
    .C(GND_0),
    .D(GND_0),
    .Z(main_basesoc_uart_tx_fifo_level0_0_mod_RNO_TMR_0)
  );
  defparam \main_basesoc_uart_tx_fifo_level0_0_mod_RNO_cZ[0]_TMR_0 .INIT = "0x4444";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55586.8-55592.2" *)
  LUT4 \main_basesoc_uart_tx_fifo_level0_0_mod_RNO_cZ[0]_TMR_1  (
    .A(sys_rst_TMR_1),
    .B(un1_main_basesoc_uart_tx_fifo_level0_TMR_1[0]),
    .C(GND_0),
    .D(GND_0),
    .Z(main_basesoc_uart_tx_fifo_level0_0_mod_RNO_TMR_1)
  );
  defparam \main_basesoc_uart_tx_fifo_level0_0_mod_RNO_cZ[0]_TMR_1 .INIT = "0x4444";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55586.8-55592.2" *)
  LUT4 \main_basesoc_uart_tx_fifo_level0_0_mod_RNO_cZ[0]_TMR_2  (
    .A(sys_rst_TMR_2),
    .B(un1_main_basesoc_uart_tx_fifo_level0_TMR_2[0]),
    .C(GND_0),
    .D(GND_0),
    .Z(main_basesoc_uart_tx_fifo_level0_0_mod_RNO_TMR_2)
  );
  defparam \main_basesoc_uart_tx_fifo_level0_0_mod_RNO_cZ[0]_TMR_2 .INIT = "0x4444";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52398.11-52404.2" *)
  FD1P3IX \main_basesoc_uart_tx_fifo_level0_mod[1]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_tx_fifo_level0_TMR_0[1]),
    .Q(un1_main_basesoc_uart_tx_fifo_level0_0_TMR_0[1]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52398.11-52404.2" *)
  FD1P3IX \main_basesoc_uart_tx_fifo_level0_mod[1]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_tx_fifo_level0_TMR_1[1]),
    .Q(un1_main_basesoc_uart_tx_fifo_level0_0_TMR_1[1]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52398.11-52404.2" *)
  FD1P3IX \main_basesoc_uart_tx_fifo_level0_mod[1]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_tx_fifo_level0_TMR_2[1]),
    .Q(un1_main_basesoc_uart_tx_fifo_level0_0_TMR_2[1]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52405.11-52411.2" *)
  FD1P3IX \main_basesoc_uart_tx_fifo_level0_mod[3]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_tx_fifo_level0_TMR_0[3]),
    .Q(un1_main_basesoc_uart_tx_fifo_level0_0_TMR_0[3]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52405.11-52411.2" *)
  FD1P3IX \main_basesoc_uart_tx_fifo_level0_mod[3]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_tx_fifo_level0_TMR_1[3]),
    .Q(un1_main_basesoc_uart_tx_fifo_level0_0_TMR_1[3]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52405.11-52411.2" *)
  FD1P3IX \main_basesoc_uart_tx_fifo_level0_mod[3]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_tx_fifo_level0_TMR_2[3]),
    .Q(un1_main_basesoc_uart_tx_fifo_level0_0_TMR_2[3]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56318.8-56324.2" *)
  LUT4 \main_basesoc_uart_tx_fifo_produce_RNO_cZ[3]_TMR_0  (
    .A(\VexRiscv.main_m1_e_0_1_TMR_0 ),
    .B(builder_csr_bankarray_csrbank3_sel_TMR_0),
    .C(main_basesoc_uart_tx_fifo_produce_TMR_0[3]),
    .D(GND_0),
    .Z(main_basesoc_uart_tx_fifo_produce_RNO_TMR_0)
  );
  defparam \main_basesoc_uart_tx_fifo_produce_RNO_cZ[3]_TMR_0 .INIT = "0x7878";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56318.8-56324.2" *)
  LUT4 \main_basesoc_uart_tx_fifo_produce_RNO_cZ[3]_TMR_1  (
    .A(\VexRiscv.main_m1_e_0_1_TMR_1 ),
    .B(builder_csr_bankarray_csrbank3_sel_TMR_1),
    .C(main_basesoc_uart_tx_fifo_produce_TMR_1[3]),
    .D(GND_0),
    .Z(main_basesoc_uart_tx_fifo_produce_RNO_TMR_1)
  );
  defparam \main_basesoc_uart_tx_fifo_produce_RNO_cZ[3]_TMR_1 .INIT = "0x7878";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56318.8-56324.2" *)
  LUT4 \main_basesoc_uart_tx_fifo_produce_RNO_cZ[3]_TMR_2  (
    .A(\VexRiscv.main_m1_e_0_1_TMR_2 ),
    .B(builder_csr_bankarray_csrbank3_sel_TMR_2),
    .C(main_basesoc_uart_tx_fifo_produce_TMR_2[3]),
    .D(GND_0),
    .Z(main_basesoc_uart_tx_fifo_produce_RNO_TMR_2)
  );
  defparam \main_basesoc_uart_tx_fifo_produce_RNO_cZ[3]_TMR_2 .INIT = "0x7878";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52370.11-52376.2" *)
  FD1P3IX \main_basesoc_uart_tx_fifo_produce_reg[0]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_tx_fifo_produce_axbxc0_TMR_0),
    .Q(main_basesoc_uart_tx_fifo_produce_TMR_0[0]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52370.11-52376.2" *)
  FD1P3IX \main_basesoc_uart_tx_fifo_produce_reg[0]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_tx_fifo_produce_axbxc0_TMR_1),
    .Q(main_basesoc_uart_tx_fifo_produce_TMR_1[0]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52370.11-52376.2" *)
  FD1P3IX \main_basesoc_uart_tx_fifo_produce_reg[0]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_tx_fifo_produce_axbxc0_TMR_2),
    .Q(main_basesoc_uart_tx_fifo_produce_TMR_2[0]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52377.11-52383.2" *)
  FD1P3IX \main_basesoc_uart_tx_fifo_produce_reg[1]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_tx_fifo_produce_axbxc1_TMR_0),
    .Q(main_basesoc_uart_tx_fifo_produce_TMR_0[1]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52377.11-52383.2" *)
  FD1P3IX \main_basesoc_uart_tx_fifo_produce_reg[1]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_tx_fifo_produce_axbxc1_TMR_1),
    .Q(main_basesoc_uart_tx_fifo_produce_TMR_1[1]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52377.11-52383.2" *)
  FD1P3IX \main_basesoc_uart_tx_fifo_produce_reg[1]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_tx_fifo_produce_axbxc1_TMR_2),
    .Q(main_basesoc_uart_tx_fifo_produce_TMR_2[1]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52384.11-52390.2" *)
  FD1P3IX \main_basesoc_uart_tx_fifo_produce_reg[2]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_tx_fifo_produce_axbxc2_TMR_0),
    .Q(main_basesoc_uart_tx_fifo_produce_TMR_0[2]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52384.11-52390.2" *)
  FD1P3IX \main_basesoc_uart_tx_fifo_produce_reg[2]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_tx_fifo_produce_axbxc2_TMR_1),
    .Q(main_basesoc_uart_tx_fifo_produce_TMR_1[2]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52384.11-52390.2" *)
  FD1P3IX \main_basesoc_uart_tx_fifo_produce_reg[2]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un1_main_basesoc_uart_tx_fifo_produce_axbxc2_TMR_2),
    .Q(main_basesoc_uart_tx_fifo_produce_TMR_2[2]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52391.11-52397.2" *)
  FD1P3IX \main_basesoc_uart_tx_fifo_produce_reg[3]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(main_basesoc_uart_tx_fifo_produce_RNO_TMR_0),
    .Q(main_basesoc_uart_tx_fifo_produce_TMR_0[3]),
    .SP(un1_main_basesoc_uart_tx_fifo_produce_axbxc3_N_13_mux_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52391.11-52397.2" *)
  FD1P3IX \main_basesoc_uart_tx_fifo_produce_reg[3]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(main_basesoc_uart_tx_fifo_produce_RNO_TMR_1),
    .Q(main_basesoc_uart_tx_fifo_produce_TMR_1[3]),
    .SP(un1_main_basesoc_uart_tx_fifo_produce_axbxc3_N_13_mux_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52391.11-52397.2" *)
  FD1P3IX \main_basesoc_uart_tx_fifo_produce_reg[3]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(main_basesoc_uart_tx_fifo_produce_RNO_TMR_2),
    .Q(main_basesoc_uart_tx_fifo_produce_TMR_2[3]),
    .SP(un1_main_basesoc_uart_tx_fifo_produce_axbxc3_N_13_mux_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52363.11-52369.2" *)
  FD1P3IX main_basesoc_uart_tx_fifo_readable_reg_TMR_0 (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(N_148_TMR_0),
    .Q(main_basesoc_uart_tx_fifo_readable_TMR_0),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52363.11-52369.2" *)
  FD1P3IX main_basesoc_uart_tx_fifo_readable_reg_TMR_1 (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(N_148_TMR_1),
    .Q(main_basesoc_uart_tx_fifo_readable_TMR_1),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52363.11-52369.2" *)
  FD1P3IX main_basesoc_uart_tx_fifo_readable_reg_TMR_2 (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(N_148_TMR_2),
    .Q(main_basesoc_uart_tx_fifo_readable_TMR_2),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52356.11-52362.2" *)
  FD1P3IX main_basesoc_uart_tx_pending_reg_TMR_0 (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(N_100_TMR_0),
    .Q(main_basesoc_uart_tx_pending_TMR_0),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52356.11-52362.2" *)
  FD1P3IX main_basesoc_uart_tx_pending_reg_TMR_1 (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(N_100_TMR_1),
    .Q(main_basesoc_uart_tx_pending_TMR_1),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52356.11-52362.2" *)
  FD1P3IX main_basesoc_uart_tx_pending_reg_TMR_2 (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(N_100_TMR_2),
    .Q(main_basesoc_uart_tx_pending_TMR_2),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52349.11-52355.2" *)
  FD1P3IX main_basesoc_uart_tx_trigger_d_reg_TMR_0 (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(un3_main_basesoc_uart_tx_fifo_syncfifo_writable_i_TMR_0),
    .Q(main_basesoc_uart_tx_trigger_d_TMR_0),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52349.11-52355.2" *)
  FD1P3IX main_basesoc_uart_tx_trigger_d_reg_TMR_1 (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(un3_main_basesoc_uart_tx_fifo_syncfifo_writable_i_TMR_1),
    .Q(main_basesoc_uart_tx_trigger_d_TMR_1),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52349.11-52355.2" *)
  FD1P3IX main_basesoc_uart_tx_trigger_d_reg_TMR_2 (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(un3_main_basesoc_uart_tx_fifo_syncfifo_writable_i_TMR_2),
    .Q(main_basesoc_uart_tx_trigger_d_TMR_2),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52342.11-52348.2" *)
  FD1P3IX main_bus_ack_reg_TMR_0 (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_bus_ack_r_0_a2_TMR_0),
    .Q(main_bus_ack_TMR_0),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52342.11-52348.2" *)
  FD1P3IX main_bus_ack_reg_TMR_1 (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_bus_ack_r_0_a2_TMR_1),
    .Q(main_bus_ack_TMR_1),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52342.11-52348.2" *)
  FD1P3IX main_bus_ack_reg_TMR_2 (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_bus_ack_r_0_a2_TMR_2),
    .Q(main_bus_ack_TMR_2),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51284.7-51287.2" *)
  INV \main_chaser_RNO[0]_TMR_0  (
    .A(main_chaser_TMR_0[13]),
    .Z(main_chaser_i_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51284.7-51287.2" *)
  INV \main_chaser_RNO[0]_TMR_1  (
    .A(main_chaser_TMR_1[13]),
    .Z(main_chaser_i_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51284.7-51287.2" *)
  INV \main_chaser_RNO[0]_TMR_2  (
    .A(main_chaser_TMR_2[13]),
    .Z(main_chaser_i_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52244.11-52250.2" *)
  FD1P3IX \main_chaser_reg[0]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(main_chaser_i_TMR_0),
    .Q(main_chaser_TMR_0[0]),
    .SP(main_done_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52244.11-52250.2" *)
  FD1P3IX \main_chaser_reg[0]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(main_chaser_i_TMR_1),
    .Q(main_chaser_TMR_1[0]),
    .SP(main_done_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52244.11-52250.2" *)
  FD1P3IX \main_chaser_reg[0]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(main_chaser_i_TMR_2),
    .Q(main_chaser_TMR_2[0]),
    .SP(main_done_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52314.11-52320.2" *)
  FD1P3IX \main_chaser_reg[10]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(main_chaser_TMR_0[9]),
    .Q(main_chaser_TMR_0[10]),
    .SP(main_done_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52314.11-52320.2" *)
  FD1P3IX \main_chaser_reg[10]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(main_chaser_TMR_1[9]),
    .Q(main_chaser_TMR_1[10]),
    .SP(main_done_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52314.11-52320.2" *)
  FD1P3IX \main_chaser_reg[10]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(main_chaser_TMR_2[9]),
    .Q(main_chaser_TMR_2[10]),
    .SP(main_done_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52321.11-52327.2" *)
  FD1P3IX \main_chaser_reg[11]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(main_chaser_TMR_0[10]),
    .Q(main_chaser_TMR_0[11]),
    .SP(main_done_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52321.11-52327.2" *)
  FD1P3IX \main_chaser_reg[11]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(main_chaser_TMR_1[10]),
    .Q(main_chaser_TMR_1[11]),
    .SP(main_done_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52321.11-52327.2" *)
  FD1P3IX \main_chaser_reg[11]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(main_chaser_TMR_2[10]),
    .Q(main_chaser_TMR_2[11]),
    .SP(main_done_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52328.11-52334.2" *)
  FD1P3IX \main_chaser_reg[12]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(main_chaser_TMR_0[11]),
    .Q(main_chaser_TMR_0[12]),
    .SP(main_done_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52328.11-52334.2" *)
  FD1P3IX \main_chaser_reg[12]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(main_chaser_TMR_1[11]),
    .Q(main_chaser_TMR_1[12]),
    .SP(main_done_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52328.11-52334.2" *)
  FD1P3IX \main_chaser_reg[12]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(main_chaser_TMR_2[11]),
    .Q(main_chaser_TMR_2[12]),
    .SP(main_done_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52335.11-52341.2" *)
  FD1P3IX \main_chaser_reg[13]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(main_chaser_TMR_0[12]),
    .Q(main_chaser_TMR_0[13]),
    .SP(main_done_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52335.11-52341.2" *)
  FD1P3IX \main_chaser_reg[13]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(main_chaser_TMR_1[12]),
    .Q(main_chaser_TMR_1[13]),
    .SP(main_done_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52335.11-52341.2" *)
  FD1P3IX \main_chaser_reg[13]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(main_chaser_TMR_2[12]),
    .Q(main_chaser_TMR_2[13]),
    .SP(main_done_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52251.11-52257.2" *)
  FD1P3IX \main_chaser_reg[1]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(main_chaser_TMR_0[0]),
    .Q(main_chaser_TMR_0[1]),
    .SP(main_done_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52251.11-52257.2" *)
  FD1P3IX \main_chaser_reg[1]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(main_chaser_TMR_1[0]),
    .Q(main_chaser_TMR_1[1]),
    .SP(main_done_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52251.11-52257.2" *)
  FD1P3IX \main_chaser_reg[1]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(main_chaser_TMR_2[0]),
    .Q(main_chaser_TMR_2[1]),
    .SP(main_done_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52258.11-52264.2" *)
  FD1P3IX \main_chaser_reg[2]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(main_chaser_TMR_0[1]),
    .Q(main_chaser_TMR_0[2]),
    .SP(main_done_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52258.11-52264.2" *)
  FD1P3IX \main_chaser_reg[2]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(main_chaser_TMR_1[1]),
    .Q(main_chaser_TMR_1[2]),
    .SP(main_done_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52258.11-52264.2" *)
  FD1P3IX \main_chaser_reg[2]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(main_chaser_TMR_2[1]),
    .Q(main_chaser_TMR_2[2]),
    .SP(main_done_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52265.11-52271.2" *)
  FD1P3IX \main_chaser_reg[3]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(main_chaser_TMR_0[2]),
    .Q(main_chaser_TMR_0[3]),
    .SP(main_done_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52265.11-52271.2" *)
  FD1P3IX \main_chaser_reg[3]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(main_chaser_TMR_1[2]),
    .Q(main_chaser_TMR_1[3]),
    .SP(main_done_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52265.11-52271.2" *)
  FD1P3IX \main_chaser_reg[3]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(main_chaser_TMR_2[2]),
    .Q(main_chaser_TMR_2[3]),
    .SP(main_done_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52272.11-52278.2" *)
  FD1P3IX \main_chaser_reg[4]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(main_chaser_TMR_0[3]),
    .Q(main_chaser_TMR_0[4]),
    .SP(main_done_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52272.11-52278.2" *)
  FD1P3IX \main_chaser_reg[4]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(main_chaser_TMR_1[3]),
    .Q(main_chaser_TMR_1[4]),
    .SP(main_done_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52272.11-52278.2" *)
  FD1P3IX \main_chaser_reg[4]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(main_chaser_TMR_2[3]),
    .Q(main_chaser_TMR_2[4]),
    .SP(main_done_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52279.11-52285.2" *)
  FD1P3IX \main_chaser_reg[5]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(main_chaser_TMR_0[4]),
    .Q(main_chaser_TMR_0[5]),
    .SP(main_done_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52279.11-52285.2" *)
  FD1P3IX \main_chaser_reg[5]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(main_chaser_TMR_1[4]),
    .Q(main_chaser_TMR_1[5]),
    .SP(main_done_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52279.11-52285.2" *)
  FD1P3IX \main_chaser_reg[5]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(main_chaser_TMR_2[4]),
    .Q(main_chaser_TMR_2[5]),
    .SP(main_done_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52286.11-52292.2" *)
  FD1P3IX \main_chaser_reg[6]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(main_chaser_TMR_0[5]),
    .Q(main_chaser_TMR_0[6]),
    .SP(main_done_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52286.11-52292.2" *)
  FD1P3IX \main_chaser_reg[6]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(main_chaser_TMR_1[5]),
    .Q(main_chaser_TMR_1[6]),
    .SP(main_done_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52286.11-52292.2" *)
  FD1P3IX \main_chaser_reg[6]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(main_chaser_TMR_2[5]),
    .Q(main_chaser_TMR_2[6]),
    .SP(main_done_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52293.11-52299.2" *)
  FD1P3IX \main_chaser_reg[7]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(main_chaser_TMR_0[6]),
    .Q(main_chaser_TMR_0[7]),
    .SP(main_done_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52293.11-52299.2" *)
  FD1P3IX \main_chaser_reg[7]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(main_chaser_TMR_1[6]),
    .Q(main_chaser_TMR_1[7]),
    .SP(main_done_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52293.11-52299.2" *)
  FD1P3IX \main_chaser_reg[7]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(main_chaser_TMR_2[6]),
    .Q(main_chaser_TMR_2[7]),
    .SP(main_done_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52300.11-52306.2" *)
  FD1P3IX \main_chaser_reg[8]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(main_chaser_TMR_0[7]),
    .Q(main_chaser_TMR_0[8]),
    .SP(main_done_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52300.11-52306.2" *)
  FD1P3IX \main_chaser_reg[8]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(main_chaser_TMR_1[7]),
    .Q(main_chaser_TMR_1[8]),
    .SP(main_done_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52300.11-52306.2" *)
  FD1P3IX \main_chaser_reg[8]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(main_chaser_TMR_2[7]),
    .Q(main_chaser_TMR_2[8]),
    .SP(main_done_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52307.11-52313.2" *)
  FD1P3IX \main_chaser_reg[9]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(main_chaser_TMR_0[8]),
    .Q(main_chaser_TMR_0[9]),
    .SP(main_done_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52307.11-52313.2" *)
  FD1P3IX \main_chaser_reg[9]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(main_chaser_TMR_1[8]),
    .Q(main_chaser_TMR_1[9]),
    .SP(main_done_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52307.11-52313.2" *)
  FD1P3IX \main_chaser_reg[9]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(main_chaser_TMR_2[8]),
    .Q(main_chaser_TMR_2[9]),
    .SP(main_done_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52090.11-52096.2" *)
  FD1P3JX \main_count[0]_TMR_0  (
    .CK(sys_clk),
    .D(main_count_RNO_TMR_0[0]),
    .PD(GND_0),
    .Q(main_count_1_TMR_0),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52090.11-52096.2" *)
  FD1P3JX \main_count[0]_TMR_1  (
    .CK(sys_clk),
    .D(main_count_RNO_TMR_1[0]),
    .PD(GND_0),
    .Q(main_count_1_TMR_1),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52090.11-52096.2" *)
  FD1P3JX \main_count[0]_TMR_2  (
    .CK(sys_clk),
    .D(main_count_RNO_TMR_2[0]),
    .PD(GND_0),
    .Q(main_count_1_TMR_2),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57929.8-57942.2" *)
  CCU2 main_count_1_cry_0_0_TMR_0 (
    .A0(VCC_TMR_0),
    .A1(main_count_1_TMR_0),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(GND_0),
    .COUT(main_count_1_cry_0_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(main_count_1_cry_0_0_S0_TMR_0),
    .S1(main_count_1_cry_0_0_S1_TMR_0)
  );
  defparam main_count_1_cry_0_0_TMR_0.INIT0 = "5033";
  defparam main_count_1_cry_0_0_TMR_0.INIT1 = "50AA";
  defparam main_count_1_cry_0_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57929.8-57942.2" *)
  CCU2 main_count_1_cry_0_0_TMR_1 (
    .A0(VCC_TMR_1),
    .A1(main_count_1_TMR_1),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(GND_0),
    .COUT(main_count_1_cry_0_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(main_count_1_cry_0_0_S0_TMR_1),
    .S1(main_count_1_cry_0_0_S1_TMR_1)
  );
  defparam main_count_1_cry_0_0_TMR_1.INIT0 = "5033";
  defparam main_count_1_cry_0_0_TMR_1.INIT1 = "50AA";
  defparam main_count_1_cry_0_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57929.8-57942.2" *)
  CCU2 main_count_1_cry_0_0_TMR_2 (
    .A0(VCC_TMR_2),
    .A1(main_count_1_TMR_2),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(GND_0),
    .COUT(main_count_1_cry_0_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(main_count_1_cry_0_0_S0_TMR_2),
    .S1(main_count_1_cry_0_0_S1_TMR_2)
  );
  defparam main_count_1_cry_0_0_TMR_2.INIT0 = "5033";
  defparam main_count_1_cry_0_0_TMR_2.INIT1 = "50AA";
  defparam main_count_1_cry_0_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57822.8-57835.2" *)
  CCU2 main_count_1_cry_11_0_TMR_0 (
    .A0(main_count_TMR_0[11]),
    .A1(main_count_TMR_0[12]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(main_count_1_cry_10_TMR_0),
    .COUT(main_count_1_cry_12_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(main_count_1_cry_11_0_S0_TMR_0),
    .S1(main_count_1_cry_11_0_S1_TMR_0)
  );
  defparam main_count_1_cry_11_0_TMR_0.INIT0 = "50AA";
  defparam main_count_1_cry_11_0_TMR_0.INIT1 = "50AA";
  defparam main_count_1_cry_11_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57822.8-57835.2" *)
  CCU2 main_count_1_cry_11_0_TMR_1 (
    .A0(main_count_TMR_1[11]),
    .A1(main_count_TMR_1[12]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(main_count_1_cry_10_TMR_1),
    .COUT(main_count_1_cry_12_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(main_count_1_cry_11_0_S0_TMR_1),
    .S1(main_count_1_cry_11_0_S1_TMR_1)
  );
  defparam main_count_1_cry_11_0_TMR_1.INIT0 = "50AA";
  defparam main_count_1_cry_11_0_TMR_1.INIT1 = "50AA";
  defparam main_count_1_cry_11_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57822.8-57835.2" *)
  CCU2 main_count_1_cry_11_0_TMR_2 (
    .A0(main_count_TMR_2[11]),
    .A1(main_count_TMR_2[12]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(main_count_1_cry_10_TMR_2),
    .COUT(main_count_1_cry_12_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(main_count_1_cry_11_0_S0_TMR_2),
    .S1(main_count_1_cry_11_0_S1_TMR_2)
  );
  defparam main_count_1_cry_11_0_TMR_2.INIT0 = "50AA";
  defparam main_count_1_cry_11_0_TMR_2.INIT1 = "50AA";
  defparam main_count_1_cry_11_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57804.8-57817.2" *)
  CCU2 main_count_1_cry_13_0_TMR_0 (
    .A0(main_count_TMR_0[13]),
    .A1(main_count_TMR_0[14]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(main_count_1_cry_12_TMR_0),
    .COUT(main_count_1_cry_14_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(main_count_1_cry_13_0_S0_TMR_0),
    .S1(main_count_1_cry_13_0_S1_TMR_0)
  );
  defparam main_count_1_cry_13_0_TMR_0.INIT0 = "50AA";
  defparam main_count_1_cry_13_0_TMR_0.INIT1 = "50AA";
  defparam main_count_1_cry_13_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57804.8-57817.2" *)
  CCU2 main_count_1_cry_13_0_TMR_1 (
    .A0(main_count_TMR_1[13]),
    .A1(main_count_TMR_1[14]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(main_count_1_cry_12_TMR_1),
    .COUT(main_count_1_cry_14_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(main_count_1_cry_13_0_S0_TMR_1),
    .S1(main_count_1_cry_13_0_S1_TMR_1)
  );
  defparam main_count_1_cry_13_0_TMR_1.INIT0 = "50AA";
  defparam main_count_1_cry_13_0_TMR_1.INIT1 = "50AA";
  defparam main_count_1_cry_13_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57804.8-57817.2" *)
  CCU2 main_count_1_cry_13_0_TMR_2 (
    .A0(main_count_TMR_2[13]),
    .A1(main_count_TMR_2[14]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(main_count_1_cry_12_TMR_2),
    .COUT(main_count_1_cry_14_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(main_count_1_cry_13_0_S0_TMR_2),
    .S1(main_count_1_cry_13_0_S1_TMR_2)
  );
  defparam main_count_1_cry_13_0_TMR_2.INIT0 = "50AA";
  defparam main_count_1_cry_13_0_TMR_2.INIT1 = "50AA";
  defparam main_count_1_cry_13_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57786.8-57799.2" *)
  CCU2 main_count_1_cry_15_0_TMR_0 (
    .A0(main_count_TMR_0[15]),
    .A1(main_count_TMR_0[16]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(main_count_1_cry_14_TMR_0),
    .COUT(main_count_1_cry_16_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(main_count_1_cry_15_0_S0_TMR_0),
    .S1(main_count_1_cry_15_0_S1_TMR_0)
  );
  defparam main_count_1_cry_15_0_TMR_0.INIT0 = "50AA";
  defparam main_count_1_cry_15_0_TMR_0.INIT1 = "50AA";
  defparam main_count_1_cry_15_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57786.8-57799.2" *)
  CCU2 main_count_1_cry_15_0_TMR_1 (
    .A0(main_count_TMR_1[15]),
    .A1(main_count_TMR_1[16]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(main_count_1_cry_14_TMR_1),
    .COUT(main_count_1_cry_16_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(main_count_1_cry_15_0_S0_TMR_1),
    .S1(main_count_1_cry_15_0_S1_TMR_1)
  );
  defparam main_count_1_cry_15_0_TMR_1.INIT0 = "50AA";
  defparam main_count_1_cry_15_0_TMR_1.INIT1 = "50AA";
  defparam main_count_1_cry_15_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57786.8-57799.2" *)
  CCU2 main_count_1_cry_15_0_TMR_2 (
    .A0(main_count_TMR_2[15]),
    .A1(main_count_TMR_2[16]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(main_count_1_cry_14_TMR_2),
    .COUT(main_count_1_cry_16_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(main_count_1_cry_15_0_S0_TMR_2),
    .S1(main_count_1_cry_15_0_S1_TMR_2)
  );
  defparam main_count_1_cry_15_0_TMR_2.INIT0 = "50AA";
  defparam main_count_1_cry_15_0_TMR_2.INIT1 = "50AA";
  defparam main_count_1_cry_15_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57768.8-57781.2" *)
  CCU2 main_count_1_cry_17_0_TMR_0 (
    .A0(main_count_TMR_0[17]),
    .A1(main_count_TMR_0[18]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(main_count_1_cry_16_TMR_0),
    .COUT(main_count_1_cry_18_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(main_count_1_cry_17_0_S0_TMR_0),
    .S1(main_count_1_cry_17_0_S1_TMR_0)
  );
  defparam main_count_1_cry_17_0_TMR_0.INIT0 = "50AA";
  defparam main_count_1_cry_17_0_TMR_0.INIT1 = "50AA";
  defparam main_count_1_cry_17_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57768.8-57781.2" *)
  CCU2 main_count_1_cry_17_0_TMR_1 (
    .A0(main_count_TMR_1[17]),
    .A1(main_count_TMR_1[18]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(main_count_1_cry_16_TMR_1),
    .COUT(main_count_1_cry_18_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(main_count_1_cry_17_0_S0_TMR_1),
    .S1(main_count_1_cry_17_0_S1_TMR_1)
  );
  defparam main_count_1_cry_17_0_TMR_1.INIT0 = "50AA";
  defparam main_count_1_cry_17_0_TMR_1.INIT1 = "50AA";
  defparam main_count_1_cry_17_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57768.8-57781.2" *)
  CCU2 main_count_1_cry_17_0_TMR_2 (
    .A0(main_count_TMR_2[17]),
    .A1(main_count_TMR_2[18]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(main_count_1_cry_16_TMR_2),
    .COUT(main_count_1_cry_18_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(main_count_1_cry_17_0_S0_TMR_2),
    .S1(main_count_1_cry_17_0_S1_TMR_2)
  );
  defparam main_count_1_cry_17_0_TMR_2.INIT0 = "50AA";
  defparam main_count_1_cry_17_0_TMR_2.INIT1 = "50AA";
  defparam main_count_1_cry_17_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57750.8-57763.2" *)
  CCU2 main_count_1_cry_19_0_TMR_0 (
    .A0(main_count_TMR_0[19]),
    .A1(main_count_TMR_0[20]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(main_count_1_cry_18_TMR_0),
    .COUT(main_count_1_cry_20_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(main_count_1_cry_19_0_S0_TMR_0),
    .S1(main_count_1_cry_19_0_S1_TMR_0)
  );
  defparam main_count_1_cry_19_0_TMR_0.INIT0 = "50AA";
  defparam main_count_1_cry_19_0_TMR_0.INIT1 = "50FF";
  defparam main_count_1_cry_19_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57750.8-57763.2" *)
  CCU2 main_count_1_cry_19_0_TMR_1 (
    .A0(main_count_TMR_1[19]),
    .A1(main_count_TMR_1[20]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(main_count_1_cry_18_TMR_1),
    .COUT(main_count_1_cry_20_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(main_count_1_cry_19_0_S0_TMR_1),
    .S1(main_count_1_cry_19_0_S1_TMR_1)
  );
  defparam main_count_1_cry_19_0_TMR_1.INIT0 = "50AA";
  defparam main_count_1_cry_19_0_TMR_1.INIT1 = "50FF";
  defparam main_count_1_cry_19_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57750.8-57763.2" *)
  CCU2 main_count_1_cry_19_0_TMR_2 (
    .A0(main_count_TMR_2[19]),
    .A1(main_count_TMR_2[20]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(main_count_1_cry_18_TMR_2),
    .COUT(main_count_1_cry_20_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(main_count_1_cry_19_0_S0_TMR_2),
    .S1(main_count_1_cry_19_0_S1_TMR_2)
  );
  defparam main_count_1_cry_19_0_TMR_2.INIT0 = "50AA";
  defparam main_count_1_cry_19_0_TMR_2.INIT1 = "50FF";
  defparam main_count_1_cry_19_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57912.8-57925.2" *)
  CCU2 main_count_1_cry_1_0_TMR_0 (
    .A0(main_count_TMR_0[1]),
    .A1(main_count_TMR_0[2]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(main_count_1_cry_0_TMR_0),
    .COUT(main_count_1_cry_2_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(main_count_1_cry_1_0_S0_TMR_0),
    .S1(main_count_1_cry_1_0_S1_TMR_0)
  );
  defparam main_count_1_cry_1_0_TMR_0.INIT0 = "50AA";
  defparam main_count_1_cry_1_0_TMR_0.INIT1 = "50AA";
  defparam main_count_1_cry_1_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57912.8-57925.2" *)
  CCU2 main_count_1_cry_1_0_TMR_1 (
    .A0(main_count_TMR_1[1]),
    .A1(main_count_TMR_1[2]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(main_count_1_cry_0_TMR_1),
    .COUT(main_count_1_cry_2_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(main_count_1_cry_1_0_S0_TMR_1),
    .S1(main_count_1_cry_1_0_S1_TMR_1)
  );
  defparam main_count_1_cry_1_0_TMR_1.INIT0 = "50AA";
  defparam main_count_1_cry_1_0_TMR_1.INIT1 = "50AA";
  defparam main_count_1_cry_1_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57912.8-57925.2" *)
  CCU2 main_count_1_cry_1_0_TMR_2 (
    .A0(main_count_TMR_2[1]),
    .A1(main_count_TMR_2[2]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(main_count_1_cry_0_TMR_2),
    .COUT(main_count_1_cry_2_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(main_count_1_cry_1_0_S0_TMR_2),
    .S1(main_count_1_cry_1_0_S1_TMR_2)
  );
  defparam main_count_1_cry_1_0_TMR_2.INIT0 = "50AA";
  defparam main_count_1_cry_1_0_TMR_2.INIT1 = "50AA";
  defparam main_count_1_cry_1_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57894.8-57907.2" *)
  CCU2 main_count_1_cry_3_0_TMR_0 (
    .A0(main_count_TMR_0[3]),
    .A1(main_count_TMR_0[4]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(main_count_1_cry_2_TMR_0),
    .COUT(main_count_1_cry_4_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(main_count_1_cry_3_0_S0_TMR_0),
    .S1(main_count_1_cry_3_0_S1_TMR_0)
  );
  defparam main_count_1_cry_3_0_TMR_0.INIT0 = "50AA";
  defparam main_count_1_cry_3_0_TMR_0.INIT1 = "50AA";
  defparam main_count_1_cry_3_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57894.8-57907.2" *)
  CCU2 main_count_1_cry_3_0_TMR_1 (
    .A0(main_count_TMR_1[3]),
    .A1(main_count_TMR_1[4]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(main_count_1_cry_2_TMR_1),
    .COUT(main_count_1_cry_4_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(main_count_1_cry_3_0_S0_TMR_1),
    .S1(main_count_1_cry_3_0_S1_TMR_1)
  );
  defparam main_count_1_cry_3_0_TMR_1.INIT0 = "50AA";
  defparam main_count_1_cry_3_0_TMR_1.INIT1 = "50AA";
  defparam main_count_1_cry_3_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57894.8-57907.2" *)
  CCU2 main_count_1_cry_3_0_TMR_2 (
    .A0(main_count_TMR_2[3]),
    .A1(main_count_TMR_2[4]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(main_count_1_cry_2_TMR_2),
    .COUT(main_count_1_cry_4_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(main_count_1_cry_3_0_S0_TMR_2),
    .S1(main_count_1_cry_3_0_S1_TMR_2)
  );
  defparam main_count_1_cry_3_0_TMR_2.INIT0 = "50AA";
  defparam main_count_1_cry_3_0_TMR_2.INIT1 = "50AA";
  defparam main_count_1_cry_3_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57876.8-57889.2" *)
  CCU2 main_count_1_cry_5_0_TMR_0 (
    .A0(main_count_TMR_0[5]),
    .A1(main_count_TMR_0[6]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(main_count_1_cry_4_TMR_0),
    .COUT(main_count_1_cry_6_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(main_count_1_cry_5_0_S0_TMR_0),
    .S1(main_count_1_cry_5_0_S1_TMR_0)
  );
  defparam main_count_1_cry_5_0_TMR_0.INIT0 = "50AA";
  defparam main_count_1_cry_5_0_TMR_0.INIT1 = "50AA";
  defparam main_count_1_cry_5_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57876.8-57889.2" *)
  CCU2 main_count_1_cry_5_0_TMR_1 (
    .A0(main_count_TMR_1[5]),
    .A1(main_count_TMR_1[6]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(main_count_1_cry_4_TMR_1),
    .COUT(main_count_1_cry_6_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(main_count_1_cry_5_0_S0_TMR_1),
    .S1(main_count_1_cry_5_0_S1_TMR_1)
  );
  defparam main_count_1_cry_5_0_TMR_1.INIT0 = "50AA";
  defparam main_count_1_cry_5_0_TMR_1.INIT1 = "50AA";
  defparam main_count_1_cry_5_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57876.8-57889.2" *)
  CCU2 main_count_1_cry_5_0_TMR_2 (
    .A0(main_count_TMR_2[5]),
    .A1(main_count_TMR_2[6]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(main_count_1_cry_4_TMR_2),
    .COUT(main_count_1_cry_6_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(main_count_1_cry_5_0_S0_TMR_2),
    .S1(main_count_1_cry_5_0_S1_TMR_2)
  );
  defparam main_count_1_cry_5_0_TMR_2.INIT0 = "50AA";
  defparam main_count_1_cry_5_0_TMR_2.INIT1 = "50AA";
  defparam main_count_1_cry_5_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57858.8-57871.2" *)
  CCU2 main_count_1_cry_7_0_TMR_0 (
    .A0(main_count_TMR_0[7]),
    .A1(main_count_TMR_0[8]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(main_count_1_cry_6_TMR_0),
    .COUT(main_count_1_cry_8_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(main_count_1_cry_7_0_S0_TMR_0),
    .S1(main_count_1_cry_7_0_S1_TMR_0)
  );
  defparam main_count_1_cry_7_0_TMR_0.INIT0 = "50AA";
  defparam main_count_1_cry_7_0_TMR_0.INIT1 = "50AA";
  defparam main_count_1_cry_7_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57858.8-57871.2" *)
  CCU2 main_count_1_cry_7_0_TMR_1 (
    .A0(main_count_TMR_1[7]),
    .A1(main_count_TMR_1[8]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(main_count_1_cry_6_TMR_1),
    .COUT(main_count_1_cry_8_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(main_count_1_cry_7_0_S0_TMR_1),
    .S1(main_count_1_cry_7_0_S1_TMR_1)
  );
  defparam main_count_1_cry_7_0_TMR_1.INIT0 = "50AA";
  defparam main_count_1_cry_7_0_TMR_1.INIT1 = "50AA";
  defparam main_count_1_cry_7_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57858.8-57871.2" *)
  CCU2 main_count_1_cry_7_0_TMR_2 (
    .A0(main_count_TMR_2[7]),
    .A1(main_count_TMR_2[8]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(main_count_1_cry_6_TMR_2),
    .COUT(main_count_1_cry_8_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(main_count_1_cry_7_0_S0_TMR_2),
    .S1(main_count_1_cry_7_0_S1_TMR_2)
  );
  defparam main_count_1_cry_7_0_TMR_2.INIT0 = "50AA";
  defparam main_count_1_cry_7_0_TMR_2.INIT1 = "50AA";
  defparam main_count_1_cry_7_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57840.8-57853.2" *)
  CCU2 main_count_1_cry_9_0_TMR_0 (
    .A0(main_count_TMR_0[9]),
    .A1(main_count_TMR_0[10]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(main_count_1_cry_8_TMR_0),
    .COUT(main_count_1_cry_10_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(main_count_1_cry_9_0_S0_TMR_0),
    .S1(main_count_1_cry_9_0_S1_TMR_0)
  );
  defparam main_count_1_cry_9_0_TMR_0.INIT0 = "50AA";
  defparam main_count_1_cry_9_0_TMR_0.INIT1 = "50AA";
  defparam main_count_1_cry_9_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57840.8-57853.2" *)
  CCU2 main_count_1_cry_9_0_TMR_1 (
    .A0(main_count_TMR_1[9]),
    .A1(main_count_TMR_1[10]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(main_count_1_cry_8_TMR_1),
    .COUT(main_count_1_cry_10_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(main_count_1_cry_9_0_S0_TMR_1),
    .S1(main_count_1_cry_9_0_S1_TMR_1)
  );
  defparam main_count_1_cry_9_0_TMR_1.INIT0 = "50AA";
  defparam main_count_1_cry_9_0_TMR_1.INIT1 = "50AA";
  defparam main_count_1_cry_9_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57840.8-57853.2" *)
  CCU2 main_count_1_cry_9_0_TMR_2 (
    .A0(main_count_TMR_2[9]),
    .A1(main_count_TMR_2[10]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(main_count_1_cry_8_TMR_2),
    .COUT(main_count_1_cry_10_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(main_count_1_cry_9_0_S0_TMR_2),
    .S1(main_count_1_cry_9_0_S1_TMR_2)
  );
  defparam main_count_1_cry_9_0_TMR_2.INIT0 = "50AA";
  defparam main_count_1_cry_9_0_TMR_2.INIT1 = "50AA";
  defparam main_count_1_cry_9_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51279.7-51282.2" *)
  INV main_count_1_s_21_0_RNO_TMR_0 (
    .A(main_count_TMR_0[21]),
    .Z(main_count_i_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51279.7-51282.2" *)
  INV main_count_1_s_21_0_RNO_TMR_1 (
    .A(main_count_TMR_1[21]),
    .Z(main_count_i_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51279.7-51282.2" *)
  INV main_count_1_s_21_0_RNO_TMR_2 (
    .A(main_count_TMR_2[21]),
    .Z(main_count_i_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57732.8-57745.2" *)
  CCU2 main_count_1_s_21_0_TMR_0 (
    .A0(main_count_i_TMR_0),
    .A1(VCC_TMR_0),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(main_count_1_cry_20_TMR_0),
    .COUT(main_count_1_s_21_0_COUT_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(main_count_1_s_21_0_S0_TMR_0),
    .S1(main_count_1_s_21_0_S1_TMR_0)
  );
  defparam main_count_1_s_21_0_TMR_0.INIT0 = "A033";
  defparam main_count_1_s_21_0_TMR_0.INIT1 = "5033";
  defparam main_count_1_s_21_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57732.8-57745.2" *)
  CCU2 main_count_1_s_21_0_TMR_1 (
    .A0(main_count_i_TMR_1),
    .A1(VCC_TMR_1),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(main_count_1_cry_20_TMR_1),
    .COUT(main_count_1_s_21_0_COUT_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(main_count_1_s_21_0_S0_TMR_1),
    .S1(main_count_1_s_21_0_S1_TMR_1)
  );
  defparam main_count_1_s_21_0_TMR_1.INIT0 = "A033";
  defparam main_count_1_s_21_0_TMR_1.INIT1 = "5033";
  defparam main_count_1_s_21_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57732.8-57745.2" *)
  CCU2 main_count_1_s_21_0_TMR_2 (
    .A0(main_count_i_TMR_2),
    .A1(VCC_TMR_2),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(main_count_1_cry_20_TMR_2),
    .COUT(main_count_1_s_21_0_COUT_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(main_count_1_s_21_0_S0_TMR_2),
    .S1(main_count_1_s_21_0_S1_TMR_2)
  );
  defparam main_count_1_s_21_0_TMR_2.INIT0 = "A033";
  defparam main_count_1_s_21_0_TMR_2.INIT1 = "5033";
  defparam main_count_1_s_21_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56074.8-56080.2" *)
  LUT4 \main_count_RNO_cZ[0]_TMR_0  (
    .A(sys_rst_TMR_0),
    .B(main_count_1_TMR_0),
    .C(GND_0),
    .D(GND_0),
    .Z(main_count_RNO_TMR_0[0])
  );
  defparam \main_count_RNO_cZ[0]_TMR_0 .INIT = "0xBBBB";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56074.8-56080.2" *)
  LUT4 \main_count_RNO_cZ[0]_TMR_1  (
    .A(sys_rst_TMR_1),
    .B(main_count_1_TMR_1),
    .C(GND_0),
    .D(GND_0),
    .Z(main_count_RNO_TMR_1[0])
  );
  defparam \main_count_RNO_cZ[0]_TMR_1 .INIT = "0xBBBB";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56074.8-56080.2" *)
  LUT4 \main_count_RNO_cZ[0]_TMR_2  (
    .A(sys_rst_TMR_2),
    .B(main_count_1_TMR_2),
    .C(GND_0),
    .D(GND_0),
    .Z(main_count_RNO_TMR_2[0])
  );
  defparam \main_count_RNO_cZ[0]_TMR_2 .INIT = "0xBBBB";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56082.8-56088.2" *)
  LUT4 \main_count_RNO_cZ[1]_TMR_0  (
    .A(sys_rst_TMR_0),
    .B(main_count_1_cry_1_0_S0_TMR_0),
    .C(GND_0),
    .D(GND_0),
    .Z(main_count_RNO_TMR_0[1])
  );
  defparam \main_count_RNO_cZ[1]_TMR_0 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56082.8-56088.2" *)
  LUT4 \main_count_RNO_cZ[1]_TMR_1  (
    .A(sys_rst_TMR_1),
    .B(main_count_1_cry_1_0_S0_TMR_1),
    .C(GND_0),
    .D(GND_0),
    .Z(main_count_RNO_TMR_1[1])
  );
  defparam \main_count_RNO_cZ[1]_TMR_1 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56082.8-56088.2" *)
  LUT4 \main_count_RNO_cZ[1]_TMR_2  (
    .A(sys_rst_TMR_2),
    .B(main_count_1_cry_1_0_S0_TMR_2),
    .C(GND_0),
    .D(GND_0),
    .Z(main_count_RNO_TMR_2[1])
  );
  defparam \main_count_RNO_cZ[1]_TMR_2 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55710.8-55716.2" *)
  LUT4 \main_count_r_0_a2_cZ[13]_TMR_0  (
    .A(sys_rst_TMR_0),
    .B(main_count_1_cry_13_0_S0_TMR_0),
    .C(main_done_TMR_0),
    .D(GND_0),
    .Z(main_count_r_0_a2_TMR_0[13])
  );
  defparam \main_count_r_0_a2_cZ[13]_TMR_0 .INIT = "0x0404";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55710.8-55716.2" *)
  LUT4 \main_count_r_0_a2_cZ[13]_TMR_1  (
    .A(sys_rst_TMR_1),
    .B(main_count_1_cry_13_0_S0_TMR_1),
    .C(main_done_TMR_1),
    .D(GND_0),
    .Z(main_count_r_0_a2_TMR_1[13])
  );
  defparam \main_count_r_0_a2_cZ[13]_TMR_1 .INIT = "0x0404";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55710.8-55716.2" *)
  LUT4 \main_count_r_0_a2_cZ[13]_TMR_2  (
    .A(sys_rst_TMR_2),
    .B(main_count_1_cry_13_0_S0_TMR_2),
    .C(main_done_TMR_2),
    .D(GND_0),
    .Z(main_count_r_0_a2_TMR_2[13])
  );
  defparam \main_count_r_0_a2_cZ[13]_TMR_2 .INIT = "0x0404";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55746.8-55752.2" *)
  LUT4 \main_count_r_0_a2_cZ[16]_TMR_0  (
    .A(sys_rst_TMR_0),
    .B(main_count_1_cry_15_0_S1_TMR_0),
    .C(main_done_TMR_0),
    .D(GND_0),
    .Z(main_count_r_0_a2_TMR_0[16])
  );
  defparam \main_count_r_0_a2_cZ[16]_TMR_0 .INIT = "0x0404";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55746.8-55752.2" *)
  LUT4 \main_count_r_0_a2_cZ[16]_TMR_1  (
    .A(sys_rst_TMR_1),
    .B(main_count_1_cry_15_0_S1_TMR_1),
    .C(main_done_TMR_1),
    .D(GND_0),
    .Z(main_count_r_0_a2_TMR_1[16])
  );
  defparam \main_count_r_0_a2_cZ[16]_TMR_1 .INIT = "0x0404";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55746.8-55752.2" *)
  LUT4 \main_count_r_0_a2_cZ[16]_TMR_2  (
    .A(sys_rst_TMR_2),
    .B(main_count_1_cry_15_0_S1_TMR_2),
    .C(main_done_TMR_2),
    .D(GND_0),
    .Z(main_count_r_0_a2_TMR_2[16])
  );
  defparam \main_count_r_0_a2_cZ[16]_TMR_2 .INIT = "0x0404";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55755.8-55761.2" *)
  LUT4 \main_count_r_0_a2_cZ[17]_TMR_0  (
    .A(sys_rst_TMR_0),
    .B(main_count_1_cry_17_0_S0_TMR_0),
    .C(main_done_TMR_0),
    .D(GND_0),
    .Z(main_count_r_0_a2_TMR_0[17])
  );
  defparam \main_count_r_0_a2_cZ[17]_TMR_0 .INIT = "0x0404";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55755.8-55761.2" *)
  LUT4 \main_count_r_0_a2_cZ[17]_TMR_1  (
    .A(sys_rst_TMR_1),
    .B(main_count_1_cry_17_0_S0_TMR_1),
    .C(main_done_TMR_1),
    .D(GND_0),
    .Z(main_count_r_0_a2_TMR_1[17])
  );
  defparam \main_count_r_0_a2_cZ[17]_TMR_1 .INIT = "0x0404";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55755.8-55761.2" *)
  LUT4 \main_count_r_0_a2_cZ[17]_TMR_2  (
    .A(sys_rst_TMR_2),
    .B(main_count_1_cry_17_0_S0_TMR_2),
    .C(main_done_TMR_2),
    .D(GND_0),
    .Z(main_count_r_0_a2_TMR_2[17])
  );
  defparam \main_count_r_0_a2_cZ[17]_TMR_2 .INIT = "0x0404";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55764.8-55770.2" *)
  LUT4 \main_count_r_0_a2_cZ[18]_TMR_0  (
    .A(sys_rst_TMR_0),
    .B(main_count_1_cry_17_0_S1_TMR_0),
    .C(main_done_TMR_0),
    .D(GND_0),
    .Z(main_count_r_0_a2_TMR_0[18])
  );
  defparam \main_count_r_0_a2_cZ[18]_TMR_0 .INIT = "0x0404";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55764.8-55770.2" *)
  LUT4 \main_count_r_0_a2_cZ[18]_TMR_1  (
    .A(sys_rst_TMR_1),
    .B(main_count_1_cry_17_0_S1_TMR_1),
    .C(main_done_TMR_1),
    .D(GND_0),
    .Z(main_count_r_0_a2_TMR_1[18])
  );
  defparam \main_count_r_0_a2_cZ[18]_TMR_1 .INIT = "0x0404";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55764.8-55770.2" *)
  LUT4 \main_count_r_0_a2_cZ[18]_TMR_2  (
    .A(sys_rst_TMR_2),
    .B(main_count_1_cry_17_0_S1_TMR_2),
    .C(main_done_TMR_2),
    .D(GND_0),
    .Z(main_count_r_0_a2_TMR_2[18])
  );
  defparam \main_count_r_0_a2_cZ[18]_TMR_2 .INIT = "0x0404";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55719.8-55725.2" *)
  LUT4 \main_count_r_0_a2_cZ[20]_TMR_0  (
    .A(sys_rst_TMR_0),
    .B(main_count_1_cry_19_0_S1_TMR_0),
    .C(main_done_TMR_0),
    .D(GND_0),
    .Z(main_count_r_0_a2_TMR_0[20])
  );
  defparam \main_count_r_0_a2_cZ[20]_TMR_0 .INIT = "0x0404";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55719.8-55725.2" *)
  LUT4 \main_count_r_0_a2_cZ[20]_TMR_1  (
    .A(sys_rst_TMR_1),
    .B(main_count_1_cry_19_0_S1_TMR_1),
    .C(main_done_TMR_1),
    .D(GND_0),
    .Z(main_count_r_0_a2_TMR_1[20])
  );
  defparam \main_count_r_0_a2_cZ[20]_TMR_1 .INIT = "0x0404";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55719.8-55725.2" *)
  LUT4 \main_count_r_0_a2_cZ[20]_TMR_2  (
    .A(sys_rst_TMR_2),
    .B(main_count_1_cry_19_0_S1_TMR_2),
    .C(main_done_TMR_2),
    .D(GND_0),
    .Z(main_count_r_0_a2_TMR_2[20])
  );
  defparam \main_count_r_0_a2_cZ[20]_TMR_2 .INIT = "0x0404";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55692.8-55698.2" *)
  LUT4 \main_count_r_0_a2_cZ[2]_TMR_0  (
    .A(sys_rst_TMR_0),
    .B(main_count_1_cry_1_0_S1_TMR_0),
    .C(main_done_TMR_0),
    .D(GND_0),
    .Z(main_count_r_0_a2_TMR_0[2])
  );
  defparam \main_count_r_0_a2_cZ[2]_TMR_0 .INIT = "0x0404";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55692.8-55698.2" *)
  LUT4 \main_count_r_0_a2_cZ[2]_TMR_1  (
    .A(sys_rst_TMR_1),
    .B(main_count_1_cry_1_0_S1_TMR_1),
    .C(main_done_TMR_1),
    .D(GND_0),
    .Z(main_count_r_0_a2_TMR_1[2])
  );
  defparam \main_count_r_0_a2_cZ[2]_TMR_1 .INIT = "0x0404";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55692.8-55698.2" *)
  LUT4 \main_count_r_0_a2_cZ[2]_TMR_2  (
    .A(sys_rst_TMR_2),
    .B(main_count_1_cry_1_0_S1_TMR_2),
    .C(main_done_TMR_2),
    .D(GND_0),
    .Z(main_count_r_0_a2_TMR_2[2])
  );
  defparam \main_count_r_0_a2_cZ[2]_TMR_2 .INIT = "0x0404";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55701.8-55707.2" *)
  LUT4 \main_count_r_0_a2_cZ[4]_TMR_0  (
    .A(sys_rst_TMR_0),
    .B(main_count_1_cry_3_0_S1_TMR_0),
    .C(main_done_TMR_0),
    .D(GND_0),
    .Z(main_count_r_0_a2_TMR_0[4])
  );
  defparam \main_count_r_0_a2_cZ[4]_TMR_0 .INIT = "0x0404";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55701.8-55707.2" *)
  LUT4 \main_count_r_0_a2_cZ[4]_TMR_1  (
    .A(sys_rst_TMR_1),
    .B(main_count_1_cry_3_0_S1_TMR_1),
    .C(main_done_TMR_1),
    .D(GND_0),
    .Z(main_count_r_0_a2_TMR_1[4])
  );
  defparam \main_count_r_0_a2_cZ[4]_TMR_1 .INIT = "0x0404";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55701.8-55707.2" *)
  LUT4 \main_count_r_0_a2_cZ[4]_TMR_2  (
    .A(sys_rst_TMR_2),
    .B(main_count_1_cry_3_0_S1_TMR_2),
    .C(main_done_TMR_2),
    .D(GND_0),
    .Z(main_count_r_0_a2_TMR_2[4])
  );
  defparam \main_count_r_0_a2_cZ[4]_TMR_2 .INIT = "0x0404";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55728.8-55734.2" *)
  LUT4 \main_count_r_0_a2_cZ[6]_TMR_0  (
    .A(sys_rst_TMR_0),
    .B(main_count_1_cry_5_0_S1_TMR_0),
    .C(main_done_TMR_0),
    .D(GND_0),
    .Z(main_count_r_0_a2_TMR_0[6])
  );
  defparam \main_count_r_0_a2_cZ[6]_TMR_0 .INIT = "0x0404";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55728.8-55734.2" *)
  LUT4 \main_count_r_0_a2_cZ[6]_TMR_1  (
    .A(sys_rst_TMR_1),
    .B(main_count_1_cry_5_0_S1_TMR_1),
    .C(main_done_TMR_1),
    .D(GND_0),
    .Z(main_count_r_0_a2_TMR_1[6])
  );
  defparam \main_count_r_0_a2_cZ[6]_TMR_1 .INIT = "0x0404";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55728.8-55734.2" *)
  LUT4 \main_count_r_0_a2_cZ[6]_TMR_2  (
    .A(sys_rst_TMR_2),
    .B(main_count_1_cry_5_0_S1_TMR_2),
    .C(main_done_TMR_2),
    .D(GND_0),
    .Z(main_count_r_0_a2_TMR_2[6])
  );
  defparam \main_count_r_0_a2_cZ[6]_TMR_2 .INIT = "0x0404";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55737.8-55743.2" *)
  LUT4 \main_count_r_0_a2_cZ[7]_TMR_0  (
    .A(sys_rst_TMR_0),
    .B(main_count_1_cry_7_0_S0_TMR_0),
    .C(main_done_TMR_0),
    .D(GND_0),
    .Z(main_count_r_0_a2_TMR_0[7])
  );
  defparam \main_count_r_0_a2_cZ[7]_TMR_0 .INIT = "0x0404";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55737.8-55743.2" *)
  LUT4 \main_count_r_0_a2_cZ[7]_TMR_1  (
    .A(sys_rst_TMR_1),
    .B(main_count_1_cry_7_0_S0_TMR_1),
    .C(main_done_TMR_1),
    .D(GND_0),
    .Z(main_count_r_0_a2_TMR_1[7])
  );
  defparam \main_count_r_0_a2_cZ[7]_TMR_1 .INIT = "0x0404";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55737.8-55743.2" *)
  LUT4 \main_count_r_0_a2_cZ[7]_TMR_2  (
    .A(sys_rst_TMR_2),
    .B(main_count_1_cry_7_0_S0_TMR_2),
    .C(main_done_TMR_2),
    .D(GND_0),
    .Z(main_count_r_0_a2_TMR_2[7])
  );
  defparam \main_count_r_0_a2_cZ[7]_TMR_2 .INIT = "0x0404";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52160.11-52166.2" *)
  FD1P3JX \main_count_reg[10]_TMR_0  (
    .CK(sys_clk),
    .D(main_count_1_cry_9_0_S1_TMR_0),
    .PD(sys_rst_TMR_0),
    .Q(main_count_TMR_0[10]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52160.11-52166.2" *)
  FD1P3JX \main_count_reg[10]_TMR_1  (
    .CK(sys_clk),
    .D(main_count_1_cry_9_0_S1_TMR_1),
    .PD(sys_rst_TMR_1),
    .Q(main_count_TMR_1[10]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52160.11-52166.2" *)
  FD1P3JX \main_count_reg[10]_TMR_2  (
    .CK(sys_clk),
    .D(main_count_1_cry_9_0_S1_TMR_2),
    .PD(sys_rst_TMR_2),
    .Q(main_count_TMR_2[10]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52167.11-52173.2" *)
  FD1P3JX \main_count_reg[11]_TMR_0  (
    .CK(sys_clk),
    .D(main_count_1_cry_11_0_S0_TMR_0),
    .PD(sys_rst_TMR_0),
    .Q(main_count_TMR_0[11]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52167.11-52173.2" *)
  FD1P3JX \main_count_reg[11]_TMR_1  (
    .CK(sys_clk),
    .D(main_count_1_cry_11_0_S0_TMR_1),
    .PD(sys_rst_TMR_1),
    .Q(main_count_TMR_1[11]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52167.11-52173.2" *)
  FD1P3JX \main_count_reg[11]_TMR_2  (
    .CK(sys_clk),
    .D(main_count_1_cry_11_0_S0_TMR_2),
    .PD(sys_rst_TMR_2),
    .Q(main_count_TMR_2[11]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52174.11-52180.2" *)
  FD1P3JX \main_count_reg[12]_TMR_0  (
    .CK(sys_clk),
    .D(main_count_1_cry_11_0_S1_TMR_0),
    .PD(sys_rst_TMR_0),
    .Q(main_count_TMR_0[12]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52174.11-52180.2" *)
  FD1P3JX \main_count_reg[12]_TMR_1  (
    .CK(sys_clk),
    .D(main_count_1_cry_11_0_S1_TMR_1),
    .PD(sys_rst_TMR_1),
    .Q(main_count_TMR_1[12]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52174.11-52180.2" *)
  FD1P3JX \main_count_reg[12]_TMR_2  (
    .CK(sys_clk),
    .D(main_count_1_cry_11_0_S1_TMR_2),
    .PD(sys_rst_TMR_2),
    .Q(main_count_TMR_2[12]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52181.11-52187.2" *)
  FD1P3IX \main_count_reg[13]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_count_r_0_a2_TMR_0[13]),
    .Q(main_count_TMR_0[13]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52181.11-52187.2" *)
  FD1P3IX \main_count_reg[13]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_count_r_0_a2_TMR_1[13]),
    .Q(main_count_TMR_1[13]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52181.11-52187.2" *)
  FD1P3IX \main_count_reg[13]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_count_r_0_a2_TMR_2[13]),
    .Q(main_count_TMR_2[13]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52188.11-52194.2" *)
  FD1P3JX \main_count_reg[14]_TMR_0  (
    .CK(sys_clk),
    .D(main_count_1_cry_13_0_S1_TMR_0),
    .PD(sys_rst_TMR_0),
    .Q(main_count_TMR_0[14]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52188.11-52194.2" *)
  FD1P3JX \main_count_reg[14]_TMR_1  (
    .CK(sys_clk),
    .D(main_count_1_cry_13_0_S1_TMR_1),
    .PD(sys_rst_TMR_1),
    .Q(main_count_TMR_1[14]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52188.11-52194.2" *)
  FD1P3JX \main_count_reg[14]_TMR_2  (
    .CK(sys_clk),
    .D(main_count_1_cry_13_0_S1_TMR_2),
    .PD(sys_rst_TMR_2),
    .Q(main_count_TMR_2[14]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52195.11-52201.2" *)
  FD1P3JX \main_count_reg[15]_TMR_0  (
    .CK(sys_clk),
    .D(main_count_1_cry_15_0_S0_TMR_0),
    .PD(sys_rst_TMR_0),
    .Q(main_count_TMR_0[15]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52195.11-52201.2" *)
  FD1P3JX \main_count_reg[15]_TMR_1  (
    .CK(sys_clk),
    .D(main_count_1_cry_15_0_S0_TMR_1),
    .PD(sys_rst_TMR_1),
    .Q(main_count_TMR_1[15]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52195.11-52201.2" *)
  FD1P3JX \main_count_reg[15]_TMR_2  (
    .CK(sys_clk),
    .D(main_count_1_cry_15_0_S0_TMR_2),
    .PD(sys_rst_TMR_2),
    .Q(main_count_TMR_2[15]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52202.11-52208.2" *)
  FD1P3IX \main_count_reg[16]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_count_r_0_a2_TMR_0[16]),
    .Q(main_count_TMR_0[16]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52202.11-52208.2" *)
  FD1P3IX \main_count_reg[16]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_count_r_0_a2_TMR_1[16]),
    .Q(main_count_TMR_1[16]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52202.11-52208.2" *)
  FD1P3IX \main_count_reg[16]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_count_r_0_a2_TMR_2[16]),
    .Q(main_count_TMR_2[16]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52209.11-52215.2" *)
  FD1P3IX \main_count_reg[17]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_count_r_0_a2_TMR_0[17]),
    .Q(main_count_TMR_0[17]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52209.11-52215.2" *)
  FD1P3IX \main_count_reg[17]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_count_r_0_a2_TMR_1[17]),
    .Q(main_count_TMR_1[17]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52209.11-52215.2" *)
  FD1P3IX \main_count_reg[17]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_count_r_0_a2_TMR_2[17]),
    .Q(main_count_TMR_2[17]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52216.11-52222.2" *)
  FD1P3IX \main_count_reg[18]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_count_r_0_a2_TMR_0[18]),
    .Q(main_count_TMR_0[18]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52216.11-52222.2" *)
  FD1P3IX \main_count_reg[18]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_count_r_0_a2_TMR_1[18]),
    .Q(main_count_TMR_1[18]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52216.11-52222.2" *)
  FD1P3IX \main_count_reg[18]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_count_r_0_a2_TMR_2[18]),
    .Q(main_count_TMR_2[18]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52223.11-52229.2" *)
  FD1P3JX \main_count_reg[19]_TMR_0  (
    .CK(sys_clk),
    .D(main_count_1_cry_19_0_S0_TMR_0),
    .PD(sys_rst_TMR_0),
    .Q(main_count_TMR_0[19]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52223.11-52229.2" *)
  FD1P3JX \main_count_reg[19]_TMR_1  (
    .CK(sys_clk),
    .D(main_count_1_cry_19_0_S0_TMR_1),
    .PD(sys_rst_TMR_1),
    .Q(main_count_TMR_1[19]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52223.11-52229.2" *)
  FD1P3JX \main_count_reg[19]_TMR_2  (
    .CK(sys_clk),
    .D(main_count_1_cry_19_0_S0_TMR_2),
    .PD(sys_rst_TMR_2),
    .Q(main_count_TMR_2[19]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52097.11-52103.2" *)
  FD1P3JX \main_count_reg[1]_TMR_0  (
    .CK(sys_clk),
    .D(main_count_RNO_TMR_0[1]),
    .PD(GND_0),
    .Q(main_count_TMR_0[1]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52097.11-52103.2" *)
  FD1P3JX \main_count_reg[1]_TMR_1  (
    .CK(sys_clk),
    .D(main_count_RNO_TMR_1[1]),
    .PD(GND_0),
    .Q(main_count_TMR_1[1]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52097.11-52103.2" *)
  FD1P3JX \main_count_reg[1]_TMR_2  (
    .CK(sys_clk),
    .D(main_count_RNO_TMR_2[1]),
    .PD(GND_0),
    .Q(main_count_TMR_2[1]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52230.11-52236.2" *)
  FD1P3IX \main_count_reg[20]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_count_r_0_a2_TMR_0[20]),
    .Q(main_count_TMR_0[20]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52230.11-52236.2" *)
  FD1P3IX \main_count_reg[20]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_count_r_0_a2_TMR_1[20]),
    .Q(main_count_TMR_1[20]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52230.11-52236.2" *)
  FD1P3IX \main_count_reg[20]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_count_r_0_a2_TMR_2[20]),
    .Q(main_count_TMR_2[20]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52237.11-52243.2" *)
  FD1P3JX \main_count_reg[21]_TMR_0  (
    .CK(sys_clk),
    .D(main_count_1_s_21_0_S0_TMR_0),
    .PD(sys_rst_TMR_0),
    .Q(main_count_TMR_0[21]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52237.11-52243.2" *)
  FD1P3JX \main_count_reg[21]_TMR_1  (
    .CK(sys_clk),
    .D(main_count_1_s_21_0_S0_TMR_1),
    .PD(sys_rst_TMR_1),
    .Q(main_count_TMR_1[21]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52237.11-52243.2" *)
  FD1P3JX \main_count_reg[21]_TMR_2  (
    .CK(sys_clk),
    .D(main_count_1_s_21_0_S0_TMR_2),
    .PD(sys_rst_TMR_2),
    .Q(main_count_TMR_2[21]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52104.11-52110.2" *)
  FD1P3IX \main_count_reg[2]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_count_r_0_a2_TMR_0[2]),
    .Q(main_count_TMR_0[2]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52104.11-52110.2" *)
  FD1P3IX \main_count_reg[2]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_count_r_0_a2_TMR_1[2]),
    .Q(main_count_TMR_1[2]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52104.11-52110.2" *)
  FD1P3IX \main_count_reg[2]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_count_r_0_a2_TMR_2[2]),
    .Q(main_count_TMR_2[2]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52111.11-52117.2" *)
  FD1P3JX \main_count_reg[3]_TMR_0  (
    .CK(sys_clk),
    .D(main_count_1_cry_3_0_S0_TMR_0),
    .PD(sys_rst_TMR_0),
    .Q(main_count_TMR_0[3]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52111.11-52117.2" *)
  FD1P3JX \main_count_reg[3]_TMR_1  (
    .CK(sys_clk),
    .D(main_count_1_cry_3_0_S0_TMR_1),
    .PD(sys_rst_TMR_1),
    .Q(main_count_TMR_1[3]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52111.11-52117.2" *)
  FD1P3JX \main_count_reg[3]_TMR_2  (
    .CK(sys_clk),
    .D(main_count_1_cry_3_0_S0_TMR_2),
    .PD(sys_rst_TMR_2),
    .Q(main_count_TMR_2[3]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52118.11-52124.2" *)
  FD1P3IX \main_count_reg[4]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_count_r_0_a2_TMR_0[4]),
    .Q(main_count_TMR_0[4]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52118.11-52124.2" *)
  FD1P3IX \main_count_reg[4]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_count_r_0_a2_TMR_1[4]),
    .Q(main_count_TMR_1[4]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52118.11-52124.2" *)
  FD1P3IX \main_count_reg[4]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_count_r_0_a2_TMR_2[4]),
    .Q(main_count_TMR_2[4]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52125.11-52131.2" *)
  FD1P3JX \main_count_reg[5]_TMR_0  (
    .CK(sys_clk),
    .D(main_count_1_cry_5_0_S0_TMR_0),
    .PD(sys_rst_TMR_0),
    .Q(main_count_TMR_0[5]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52125.11-52131.2" *)
  FD1P3JX \main_count_reg[5]_TMR_1  (
    .CK(sys_clk),
    .D(main_count_1_cry_5_0_S0_TMR_1),
    .PD(sys_rst_TMR_1),
    .Q(main_count_TMR_1[5]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52125.11-52131.2" *)
  FD1P3JX \main_count_reg[5]_TMR_2  (
    .CK(sys_clk),
    .D(main_count_1_cry_5_0_S0_TMR_2),
    .PD(sys_rst_TMR_2),
    .Q(main_count_TMR_2[5]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52132.11-52138.2" *)
  FD1P3IX \main_count_reg[6]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_count_r_0_a2_TMR_0[6]),
    .Q(main_count_TMR_0[6]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52132.11-52138.2" *)
  FD1P3IX \main_count_reg[6]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_count_r_0_a2_TMR_1[6]),
    .Q(main_count_TMR_1[6]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52132.11-52138.2" *)
  FD1P3IX \main_count_reg[6]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_count_r_0_a2_TMR_2[6]),
    .Q(main_count_TMR_2[6]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52139.11-52145.2" *)
  FD1P3IX \main_count_reg[7]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_count_r_0_a2_TMR_0[7]),
    .Q(main_count_TMR_0[7]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52139.11-52145.2" *)
  FD1P3IX \main_count_reg[7]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_count_r_0_a2_TMR_1[7]),
    .Q(main_count_TMR_1[7]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52139.11-52145.2" *)
  FD1P3IX \main_count_reg[7]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_count_r_0_a2_TMR_2[7]),
    .Q(main_count_TMR_2[7]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52146.11-52152.2" *)
  FD1P3JX \main_count_reg[8]_TMR_0  (
    .CK(sys_clk),
    .D(main_count_1_cry_7_0_S1_TMR_0),
    .PD(sys_rst_TMR_0),
    .Q(main_count_TMR_0[8]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52146.11-52152.2" *)
  FD1P3JX \main_count_reg[8]_TMR_1  (
    .CK(sys_clk),
    .D(main_count_1_cry_7_0_S1_TMR_1),
    .PD(sys_rst_TMR_1),
    .Q(main_count_TMR_1[8]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52146.11-52152.2" *)
  FD1P3JX \main_count_reg[8]_TMR_2  (
    .CK(sys_clk),
    .D(main_count_1_cry_7_0_S1_TMR_2),
    .PD(sys_rst_TMR_2),
    .Q(main_count_TMR_2[8]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52153.11-52159.2" *)
  FD1P3JX \main_count_reg[9]_TMR_0  (
    .CK(sys_clk),
    .D(main_count_1_cry_9_0_S0_TMR_0),
    .PD(sys_rst_TMR_0),
    .Q(main_count_TMR_0[9]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52153.11-52159.2" *)
  FD1P3JX \main_count_reg[9]_TMR_1  (
    .CK(sys_clk),
    .D(main_count_1_cry_9_0_S0_TMR_1),
    .PD(sys_rst_TMR_1),
    .Q(main_count_TMR_1[9]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52153.11-52159.2" *)
  FD1P3JX \main_count_reg[9]_TMR_2  (
    .CK(sys_clk),
    .D(main_count_1_cry_9_0_S0_TMR_2),
    .PD(sys_rst_TMR_2),
    .Q(main_count_TMR_2[9]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55808.8-55814.2" *)
  LUT4 \main_crg_por_count_RNO_cZ[0]_TMR_0  (
    .A(por_rst_TMR_0),
    .B(main_crg_por_count_TMR_0[0]),
    .C(main_crg_por_done_12_TMR_0),
    .D(main_crg_por_done_13_TMR_0),
    .Z(main_crg_por_count_RNO_TMR_0[0])
  );
  defparam \main_crg_por_count_RNO_cZ[0]_TMR_0 .INIT = "0xEBBB";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55808.8-55814.2" *)
  LUT4 \main_crg_por_count_RNO_cZ[0]_TMR_1  (
    .A(por_rst_TMR_1),
    .B(main_crg_por_count_TMR_1[0]),
    .C(main_crg_por_done_12_TMR_1),
    .D(main_crg_por_done_13_TMR_1),
    .Z(main_crg_por_count_RNO_TMR_1[0])
  );
  defparam \main_crg_por_count_RNO_cZ[0]_TMR_1 .INIT = "0xEBBB";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55808.8-55814.2" *)
  LUT4 \main_crg_por_count_RNO_cZ[0]_TMR_2  (
    .A(por_rst_TMR_2),
    .B(main_crg_por_count_TMR_2[0]),
    .C(main_crg_por_done_12_TMR_2),
    .D(main_crg_por_done_13_TMR_2),
    .Z(main_crg_por_count_RNO_TMR_2[0])
  );
  defparam \main_crg_por_count_RNO_cZ[0]_TMR_2 .INIT = "0xEBBB";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56162.8-56168.2" *)
  LUT4 \main_crg_por_count_RNO_cZ[10]_TMR_0  (
    .A(por_rst_TMR_0),
    .B(un1_main_crg_por_count_cry_9_0_S1_TMR_0),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_count_RNO_TMR_0[10])
  );
  defparam \main_crg_por_count_RNO_cZ[10]_TMR_0 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56162.8-56168.2" *)
  LUT4 \main_crg_por_count_RNO_cZ[10]_TMR_1  (
    .A(por_rst_TMR_1),
    .B(un1_main_crg_por_count_cry_9_0_S1_TMR_1),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_count_RNO_TMR_1[10])
  );
  defparam \main_crg_por_count_RNO_cZ[10]_TMR_1 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56162.8-56168.2" *)
  LUT4 \main_crg_por_count_RNO_cZ[10]_TMR_2  (
    .A(por_rst_TMR_2),
    .B(un1_main_crg_por_count_cry_9_0_S1_TMR_2),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_count_RNO_TMR_2[10])
  );
  defparam \main_crg_por_count_RNO_cZ[10]_TMR_2 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56170.8-56176.2" *)
  LUT4 \main_crg_por_count_RNO_cZ[11]_TMR_0  (
    .A(por_rst_TMR_0),
    .B(un1_main_crg_por_count_cry_11_0_S0_TMR_0),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_count_RNO_TMR_0[11])
  );
  defparam \main_crg_por_count_RNO_cZ[11]_TMR_0 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56170.8-56176.2" *)
  LUT4 \main_crg_por_count_RNO_cZ[11]_TMR_1  (
    .A(por_rst_TMR_1),
    .B(un1_main_crg_por_count_cry_11_0_S0_TMR_1),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_count_RNO_TMR_1[11])
  );
  defparam \main_crg_por_count_RNO_cZ[11]_TMR_1 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56170.8-56176.2" *)
  LUT4 \main_crg_por_count_RNO_cZ[11]_TMR_2  (
    .A(por_rst_TMR_2),
    .B(un1_main_crg_por_count_cry_11_0_S0_TMR_2),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_count_RNO_TMR_2[11])
  );
  defparam \main_crg_por_count_RNO_cZ[11]_TMR_2 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56178.8-56184.2" *)
  LUT4 \main_crg_por_count_RNO_cZ[12]_TMR_0  (
    .A(por_rst_TMR_0),
    .B(un1_main_crg_por_count_cry_11_0_S1_TMR_0),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_count_RNO_TMR_0[12])
  );
  defparam \main_crg_por_count_RNO_cZ[12]_TMR_0 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56178.8-56184.2" *)
  LUT4 \main_crg_por_count_RNO_cZ[12]_TMR_1  (
    .A(por_rst_TMR_1),
    .B(un1_main_crg_por_count_cry_11_0_S1_TMR_1),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_count_RNO_TMR_1[12])
  );
  defparam \main_crg_por_count_RNO_cZ[12]_TMR_1 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56178.8-56184.2" *)
  LUT4 \main_crg_por_count_RNO_cZ[12]_TMR_2  (
    .A(por_rst_TMR_2),
    .B(un1_main_crg_por_count_cry_11_0_S1_TMR_2),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_count_RNO_TMR_2[12])
  );
  defparam \main_crg_por_count_RNO_cZ[12]_TMR_2 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56186.8-56192.2" *)
  LUT4 \main_crg_por_count_RNO_cZ[13]_TMR_0  (
    .A(por_rst_TMR_0),
    .B(un1_main_crg_por_count_cry_13_0_S0_TMR_0),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_count_RNO_TMR_0[13])
  );
  defparam \main_crg_por_count_RNO_cZ[13]_TMR_0 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56186.8-56192.2" *)
  LUT4 \main_crg_por_count_RNO_cZ[13]_TMR_1  (
    .A(por_rst_TMR_1),
    .B(un1_main_crg_por_count_cry_13_0_S0_TMR_1),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_count_RNO_TMR_1[13])
  );
  defparam \main_crg_por_count_RNO_cZ[13]_TMR_1 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56186.8-56192.2" *)
  LUT4 \main_crg_por_count_RNO_cZ[13]_TMR_2  (
    .A(por_rst_TMR_2),
    .B(un1_main_crg_por_count_cry_13_0_S0_TMR_2),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_count_RNO_TMR_2[13])
  );
  defparam \main_crg_por_count_RNO_cZ[13]_TMR_2 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56194.8-56200.2" *)
  LUT4 \main_crg_por_count_RNO_cZ[14]_TMR_0  (
    .A(por_rst_TMR_0),
    .B(un1_main_crg_por_count_cry_13_0_S1_TMR_0),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_count_RNO_TMR_0[14])
  );
  defparam \main_crg_por_count_RNO_cZ[14]_TMR_0 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56194.8-56200.2" *)
  LUT4 \main_crg_por_count_RNO_cZ[14]_TMR_1  (
    .A(por_rst_TMR_1),
    .B(un1_main_crg_por_count_cry_13_0_S1_TMR_1),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_count_RNO_TMR_1[14])
  );
  defparam \main_crg_por_count_RNO_cZ[14]_TMR_1 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56194.8-56200.2" *)
  LUT4 \main_crg_por_count_RNO_cZ[14]_TMR_2  (
    .A(por_rst_TMR_2),
    .B(un1_main_crg_por_count_cry_13_0_S1_TMR_2),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_count_RNO_TMR_2[14])
  );
  defparam \main_crg_por_count_RNO_cZ[14]_TMR_2 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56202.8-56208.2" *)
  LUT4 \main_crg_por_count_RNO_cZ[15]_TMR_0  (
    .A(por_rst_TMR_0),
    .B(un1_main_crg_por_count_s_15_0_S0_TMR_0),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_count_RNO_TMR_0[15])
  );
  defparam \main_crg_por_count_RNO_cZ[15]_TMR_0 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56202.8-56208.2" *)
  LUT4 \main_crg_por_count_RNO_cZ[15]_TMR_1  (
    .A(por_rst_TMR_1),
    .B(un1_main_crg_por_count_s_15_0_S0_TMR_1),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_count_RNO_TMR_1[15])
  );
  defparam \main_crg_por_count_RNO_cZ[15]_TMR_1 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56202.8-56208.2" *)
  LUT4 \main_crg_por_count_RNO_cZ[15]_TMR_2  (
    .A(por_rst_TMR_2),
    .B(un1_main_crg_por_count_s_15_0_S0_TMR_2),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_count_RNO_TMR_2[15])
  );
  defparam \main_crg_por_count_RNO_cZ[15]_TMR_2 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56090.8-56096.2" *)
  LUT4 \main_crg_por_count_RNO_cZ[1]_TMR_0  (
    .A(por_rst_TMR_0),
    .B(un1_main_crg_por_count_cry_1_0_S0_TMR_0),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_count_RNO_TMR_0[1])
  );
  defparam \main_crg_por_count_RNO_cZ[1]_TMR_0 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56090.8-56096.2" *)
  LUT4 \main_crg_por_count_RNO_cZ[1]_TMR_1  (
    .A(por_rst_TMR_1),
    .B(un1_main_crg_por_count_cry_1_0_S0_TMR_1),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_count_RNO_TMR_1[1])
  );
  defparam \main_crg_por_count_RNO_cZ[1]_TMR_1 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56090.8-56096.2" *)
  LUT4 \main_crg_por_count_RNO_cZ[1]_TMR_2  (
    .A(por_rst_TMR_2),
    .B(un1_main_crg_por_count_cry_1_0_S0_TMR_2),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_count_RNO_TMR_2[1])
  );
  defparam \main_crg_por_count_RNO_cZ[1]_TMR_2 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56098.8-56104.2" *)
  LUT4 \main_crg_por_count_RNO_cZ[2]_TMR_0  (
    .A(por_rst_TMR_0),
    .B(un1_main_crg_por_count_cry_1_0_S1_TMR_0),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_count_RNO_TMR_0[2])
  );
  defparam \main_crg_por_count_RNO_cZ[2]_TMR_0 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56098.8-56104.2" *)
  LUT4 \main_crg_por_count_RNO_cZ[2]_TMR_1  (
    .A(por_rst_TMR_1),
    .B(un1_main_crg_por_count_cry_1_0_S1_TMR_1),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_count_RNO_TMR_1[2])
  );
  defparam \main_crg_por_count_RNO_cZ[2]_TMR_1 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56098.8-56104.2" *)
  LUT4 \main_crg_por_count_RNO_cZ[2]_TMR_2  (
    .A(por_rst_TMR_2),
    .B(un1_main_crg_por_count_cry_1_0_S1_TMR_2),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_count_RNO_TMR_2[2])
  );
  defparam \main_crg_por_count_RNO_cZ[2]_TMR_2 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56106.8-56112.2" *)
  LUT4 \main_crg_por_count_RNO_cZ[3]_TMR_0  (
    .A(por_rst_TMR_0),
    .B(un1_main_crg_por_count_cry_3_0_S0_TMR_0),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_count_RNO_TMR_0[3])
  );
  defparam \main_crg_por_count_RNO_cZ[3]_TMR_0 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56106.8-56112.2" *)
  LUT4 \main_crg_por_count_RNO_cZ[3]_TMR_1  (
    .A(por_rst_TMR_1),
    .B(un1_main_crg_por_count_cry_3_0_S0_TMR_1),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_count_RNO_TMR_1[3])
  );
  defparam \main_crg_por_count_RNO_cZ[3]_TMR_1 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56106.8-56112.2" *)
  LUT4 \main_crg_por_count_RNO_cZ[3]_TMR_2  (
    .A(por_rst_TMR_2),
    .B(un1_main_crg_por_count_cry_3_0_S0_TMR_2),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_count_RNO_TMR_2[3])
  );
  defparam \main_crg_por_count_RNO_cZ[3]_TMR_2 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56114.8-56120.2" *)
  LUT4 \main_crg_por_count_RNO_cZ[4]_TMR_0  (
    .A(por_rst_TMR_0),
    .B(un1_main_crg_por_count_cry_3_0_S1_TMR_0),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_count_RNO_TMR_0[4])
  );
  defparam \main_crg_por_count_RNO_cZ[4]_TMR_0 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56114.8-56120.2" *)
  LUT4 \main_crg_por_count_RNO_cZ[4]_TMR_1  (
    .A(por_rst_TMR_1),
    .B(un1_main_crg_por_count_cry_3_0_S1_TMR_1),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_count_RNO_TMR_1[4])
  );
  defparam \main_crg_por_count_RNO_cZ[4]_TMR_1 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56114.8-56120.2" *)
  LUT4 \main_crg_por_count_RNO_cZ[4]_TMR_2  (
    .A(por_rst_TMR_2),
    .B(un1_main_crg_por_count_cry_3_0_S1_TMR_2),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_count_RNO_TMR_2[4])
  );
  defparam \main_crg_por_count_RNO_cZ[4]_TMR_2 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56122.8-56128.2" *)
  LUT4 \main_crg_por_count_RNO_cZ[5]_TMR_0  (
    .A(por_rst_TMR_0),
    .B(un1_main_crg_por_count_cry_5_0_S0_TMR_0),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_count_RNO_TMR_0[5])
  );
  defparam \main_crg_por_count_RNO_cZ[5]_TMR_0 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56122.8-56128.2" *)
  LUT4 \main_crg_por_count_RNO_cZ[5]_TMR_1  (
    .A(por_rst_TMR_1),
    .B(un1_main_crg_por_count_cry_5_0_S0_TMR_1),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_count_RNO_TMR_1[5])
  );
  defparam \main_crg_por_count_RNO_cZ[5]_TMR_1 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56122.8-56128.2" *)
  LUT4 \main_crg_por_count_RNO_cZ[5]_TMR_2  (
    .A(por_rst_TMR_2),
    .B(un1_main_crg_por_count_cry_5_0_S0_TMR_2),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_count_RNO_TMR_2[5])
  );
  defparam \main_crg_por_count_RNO_cZ[5]_TMR_2 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56130.8-56136.2" *)
  LUT4 \main_crg_por_count_RNO_cZ[6]_TMR_0  (
    .A(por_rst_TMR_0),
    .B(un1_main_crg_por_count_cry_5_0_S1_TMR_0),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_count_RNO_TMR_0[6])
  );
  defparam \main_crg_por_count_RNO_cZ[6]_TMR_0 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56130.8-56136.2" *)
  LUT4 \main_crg_por_count_RNO_cZ[6]_TMR_1  (
    .A(por_rst_TMR_1),
    .B(un1_main_crg_por_count_cry_5_0_S1_TMR_1),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_count_RNO_TMR_1[6])
  );
  defparam \main_crg_por_count_RNO_cZ[6]_TMR_1 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56130.8-56136.2" *)
  LUT4 \main_crg_por_count_RNO_cZ[6]_TMR_2  (
    .A(por_rst_TMR_2),
    .B(un1_main_crg_por_count_cry_5_0_S1_TMR_2),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_count_RNO_TMR_2[6])
  );
  defparam \main_crg_por_count_RNO_cZ[6]_TMR_2 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56138.8-56144.2" *)
  LUT4 \main_crg_por_count_RNO_cZ[7]_TMR_0  (
    .A(por_rst_TMR_0),
    .B(un1_main_crg_por_count_cry_7_0_S0_TMR_0),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_count_RNO_TMR_0[7])
  );
  defparam \main_crg_por_count_RNO_cZ[7]_TMR_0 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56138.8-56144.2" *)
  LUT4 \main_crg_por_count_RNO_cZ[7]_TMR_1  (
    .A(por_rst_TMR_1),
    .B(un1_main_crg_por_count_cry_7_0_S0_TMR_1),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_count_RNO_TMR_1[7])
  );
  defparam \main_crg_por_count_RNO_cZ[7]_TMR_1 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56138.8-56144.2" *)
  LUT4 \main_crg_por_count_RNO_cZ[7]_TMR_2  (
    .A(por_rst_TMR_2),
    .B(un1_main_crg_por_count_cry_7_0_S0_TMR_2),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_count_RNO_TMR_2[7])
  );
  defparam \main_crg_por_count_RNO_cZ[7]_TMR_2 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56146.8-56152.2" *)
  LUT4 \main_crg_por_count_RNO_cZ[8]_TMR_0  (
    .A(por_rst_TMR_0),
    .B(un1_main_crg_por_count_cry_7_0_S1_TMR_0),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_count_RNO_TMR_0[8])
  );
  defparam \main_crg_por_count_RNO_cZ[8]_TMR_0 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56146.8-56152.2" *)
  LUT4 \main_crg_por_count_RNO_cZ[8]_TMR_1  (
    .A(por_rst_TMR_1),
    .B(un1_main_crg_por_count_cry_7_0_S1_TMR_1),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_count_RNO_TMR_1[8])
  );
  defparam \main_crg_por_count_RNO_cZ[8]_TMR_1 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56146.8-56152.2" *)
  LUT4 \main_crg_por_count_RNO_cZ[8]_TMR_2  (
    .A(por_rst_TMR_2),
    .B(un1_main_crg_por_count_cry_7_0_S1_TMR_2),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_count_RNO_TMR_2[8])
  );
  defparam \main_crg_por_count_RNO_cZ[8]_TMR_2 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56154.8-56160.2" *)
  LUT4 \main_crg_por_count_RNO_cZ[9]_TMR_0  (
    .A(por_rst_TMR_0),
    .B(un1_main_crg_por_count_cry_9_0_S0_TMR_0),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_count_RNO_TMR_0[9])
  );
  defparam \main_crg_por_count_RNO_cZ[9]_TMR_0 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56154.8-56160.2" *)
  LUT4 \main_crg_por_count_RNO_cZ[9]_TMR_1  (
    .A(por_rst_TMR_1),
    .B(un1_main_crg_por_count_cry_9_0_S0_TMR_1),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_count_RNO_TMR_1[9])
  );
  defparam \main_crg_por_count_RNO_cZ[9]_TMR_1 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56154.8-56160.2" *)
  LUT4 \main_crg_por_count_RNO_cZ[9]_TMR_2  (
    .A(por_rst_TMR_2),
    .B(un1_main_crg_por_count_cry_9_0_S0_TMR_2),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_count_RNO_TMR_2[9])
  );
  defparam \main_crg_por_count_RNO_cZ[9]_TMR_2 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51978.11-51984.2" *)
  FD1P3JX \main_crg_por_count_reg[0]_TMR_0  (
    .CK(main_crg_clkout),
    .D(main_crg_por_count_RNO_TMR_0[0]),
    .PD(GND_0),
    .Q(main_crg_por_count_TMR_0[0]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51978.11-51984.2" *)
  FD1P3JX \main_crg_por_count_reg[0]_TMR_1  (
    .CK(main_crg_clkout),
    .D(main_crg_por_count_RNO_TMR_1[0]),
    .PD(GND_0),
    .Q(main_crg_por_count_TMR_1[0]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51978.11-51984.2" *)
  FD1P3JX \main_crg_por_count_reg[0]_TMR_2  (
    .CK(main_crg_clkout),
    .D(main_crg_por_count_RNO_TMR_2[0]),
    .PD(GND_0),
    .Q(main_crg_por_count_TMR_2[0]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52048.11-52054.2" *)
  FD1P3JX \main_crg_por_count_reg[10]_TMR_0  (
    .CK(main_crg_clkout),
    .D(main_crg_por_count_RNO_TMR_0[10]),
    .PD(GND_0),
    .Q(main_crg_por_count_TMR_0[10]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52048.11-52054.2" *)
  FD1P3JX \main_crg_por_count_reg[10]_TMR_1  (
    .CK(main_crg_clkout),
    .D(main_crg_por_count_RNO_TMR_1[10]),
    .PD(GND_0),
    .Q(main_crg_por_count_TMR_1[10]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52048.11-52054.2" *)
  FD1P3JX \main_crg_por_count_reg[10]_TMR_2  (
    .CK(main_crg_clkout),
    .D(main_crg_por_count_RNO_TMR_2[10]),
    .PD(GND_0),
    .Q(main_crg_por_count_TMR_2[10]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52055.11-52061.2" *)
  FD1P3JX \main_crg_por_count_reg[11]_TMR_0  (
    .CK(main_crg_clkout),
    .D(main_crg_por_count_RNO_TMR_0[11]),
    .PD(GND_0),
    .Q(main_crg_por_count_TMR_0[11]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52055.11-52061.2" *)
  FD1P3JX \main_crg_por_count_reg[11]_TMR_1  (
    .CK(main_crg_clkout),
    .D(main_crg_por_count_RNO_TMR_1[11]),
    .PD(GND_0),
    .Q(main_crg_por_count_TMR_1[11]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52055.11-52061.2" *)
  FD1P3JX \main_crg_por_count_reg[11]_TMR_2  (
    .CK(main_crg_clkout),
    .D(main_crg_por_count_RNO_TMR_2[11]),
    .PD(GND_0),
    .Q(main_crg_por_count_TMR_2[11]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52062.11-52068.2" *)
  FD1P3JX \main_crg_por_count_reg[12]_TMR_0  (
    .CK(main_crg_clkout),
    .D(main_crg_por_count_RNO_TMR_0[12]),
    .PD(GND_0),
    .Q(main_crg_por_count_TMR_0[12]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52062.11-52068.2" *)
  FD1P3JX \main_crg_por_count_reg[12]_TMR_1  (
    .CK(main_crg_clkout),
    .D(main_crg_por_count_RNO_TMR_1[12]),
    .PD(GND_0),
    .Q(main_crg_por_count_TMR_1[12]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52062.11-52068.2" *)
  FD1P3JX \main_crg_por_count_reg[12]_TMR_2  (
    .CK(main_crg_clkout),
    .D(main_crg_por_count_RNO_TMR_2[12]),
    .PD(GND_0),
    .Q(main_crg_por_count_TMR_2[12]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52069.11-52075.2" *)
  FD1P3JX \main_crg_por_count_reg[13]_TMR_0  (
    .CK(main_crg_clkout),
    .D(main_crg_por_count_RNO_TMR_0[13]),
    .PD(GND_0),
    .Q(main_crg_por_count_TMR_0[13]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52069.11-52075.2" *)
  FD1P3JX \main_crg_por_count_reg[13]_TMR_1  (
    .CK(main_crg_clkout),
    .D(main_crg_por_count_RNO_TMR_1[13]),
    .PD(GND_0),
    .Q(main_crg_por_count_TMR_1[13]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52069.11-52075.2" *)
  FD1P3JX \main_crg_por_count_reg[13]_TMR_2  (
    .CK(main_crg_clkout),
    .D(main_crg_por_count_RNO_TMR_2[13]),
    .PD(GND_0),
    .Q(main_crg_por_count_TMR_2[13]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52076.11-52082.2" *)
  FD1P3JX \main_crg_por_count_reg[14]_TMR_0  (
    .CK(main_crg_clkout),
    .D(main_crg_por_count_RNO_TMR_0[14]),
    .PD(GND_0),
    .Q(main_crg_por_count_TMR_0[14]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52076.11-52082.2" *)
  FD1P3JX \main_crg_por_count_reg[14]_TMR_1  (
    .CK(main_crg_clkout),
    .D(main_crg_por_count_RNO_TMR_1[14]),
    .PD(GND_0),
    .Q(main_crg_por_count_TMR_1[14]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52076.11-52082.2" *)
  FD1P3JX \main_crg_por_count_reg[14]_TMR_2  (
    .CK(main_crg_clkout),
    .D(main_crg_por_count_RNO_TMR_2[14]),
    .PD(GND_0),
    .Q(main_crg_por_count_TMR_2[14]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52083.11-52089.2" *)
  FD1P3JX \main_crg_por_count_reg[15]_TMR_0  (
    .CK(main_crg_clkout),
    .D(main_crg_por_count_RNO_TMR_0[15]),
    .PD(GND_0),
    .Q(main_crg_por_count_TMR_0[15]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52083.11-52089.2" *)
  FD1P3JX \main_crg_por_count_reg[15]_TMR_1  (
    .CK(main_crg_clkout),
    .D(main_crg_por_count_RNO_TMR_1[15]),
    .PD(GND_0),
    .Q(main_crg_por_count_TMR_1[15]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52083.11-52089.2" *)
  FD1P3JX \main_crg_por_count_reg[15]_TMR_2  (
    .CK(main_crg_clkout),
    .D(main_crg_por_count_RNO_TMR_2[15]),
    .PD(GND_0),
    .Q(main_crg_por_count_TMR_2[15]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51985.11-51991.2" *)
  FD1P3JX \main_crg_por_count_reg[1]_TMR_0  (
    .CK(main_crg_clkout),
    .D(main_crg_por_count_RNO_TMR_0[1]),
    .PD(GND_0),
    .Q(main_crg_por_count_TMR_0[1]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51985.11-51991.2" *)
  FD1P3JX \main_crg_por_count_reg[1]_TMR_1  (
    .CK(main_crg_clkout),
    .D(main_crg_por_count_RNO_TMR_1[1]),
    .PD(GND_0),
    .Q(main_crg_por_count_TMR_1[1]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51985.11-51991.2" *)
  FD1P3JX \main_crg_por_count_reg[1]_TMR_2  (
    .CK(main_crg_clkout),
    .D(main_crg_por_count_RNO_TMR_2[1]),
    .PD(GND_0),
    .Q(main_crg_por_count_TMR_2[1]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51992.11-51998.2" *)
  FD1P3JX \main_crg_por_count_reg[2]_TMR_0  (
    .CK(main_crg_clkout),
    .D(main_crg_por_count_RNO_TMR_0[2]),
    .PD(GND_0),
    .Q(main_crg_por_count_TMR_0[2]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51992.11-51998.2" *)
  FD1P3JX \main_crg_por_count_reg[2]_TMR_1  (
    .CK(main_crg_clkout),
    .D(main_crg_por_count_RNO_TMR_1[2]),
    .PD(GND_0),
    .Q(main_crg_por_count_TMR_1[2]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51992.11-51998.2" *)
  FD1P3JX \main_crg_por_count_reg[2]_TMR_2  (
    .CK(main_crg_clkout),
    .D(main_crg_por_count_RNO_TMR_2[2]),
    .PD(GND_0),
    .Q(main_crg_por_count_TMR_2[2]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51999.11-52005.2" *)
  FD1P3JX \main_crg_por_count_reg[3]_TMR_0  (
    .CK(main_crg_clkout),
    .D(main_crg_por_count_RNO_TMR_0[3]),
    .PD(GND_0),
    .Q(main_crg_por_count_TMR_0[3]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51999.11-52005.2" *)
  FD1P3JX \main_crg_por_count_reg[3]_TMR_1  (
    .CK(main_crg_clkout),
    .D(main_crg_por_count_RNO_TMR_1[3]),
    .PD(GND_0),
    .Q(main_crg_por_count_TMR_1[3]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51999.11-52005.2" *)
  FD1P3JX \main_crg_por_count_reg[3]_TMR_2  (
    .CK(main_crg_clkout),
    .D(main_crg_por_count_RNO_TMR_2[3]),
    .PD(GND_0),
    .Q(main_crg_por_count_TMR_2[3]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52006.11-52012.2" *)
  FD1P3JX \main_crg_por_count_reg[4]_TMR_0  (
    .CK(main_crg_clkout),
    .D(main_crg_por_count_RNO_TMR_0[4]),
    .PD(GND_0),
    .Q(main_crg_por_count_TMR_0[4]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52006.11-52012.2" *)
  FD1P3JX \main_crg_por_count_reg[4]_TMR_1  (
    .CK(main_crg_clkout),
    .D(main_crg_por_count_RNO_TMR_1[4]),
    .PD(GND_0),
    .Q(main_crg_por_count_TMR_1[4]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52006.11-52012.2" *)
  FD1P3JX \main_crg_por_count_reg[4]_TMR_2  (
    .CK(main_crg_clkout),
    .D(main_crg_por_count_RNO_TMR_2[4]),
    .PD(GND_0),
    .Q(main_crg_por_count_TMR_2[4]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52013.11-52019.2" *)
  FD1P3JX \main_crg_por_count_reg[5]_TMR_0  (
    .CK(main_crg_clkout),
    .D(main_crg_por_count_RNO_TMR_0[5]),
    .PD(GND_0),
    .Q(main_crg_por_count_TMR_0[5]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52013.11-52019.2" *)
  FD1P3JX \main_crg_por_count_reg[5]_TMR_1  (
    .CK(main_crg_clkout),
    .D(main_crg_por_count_RNO_TMR_1[5]),
    .PD(GND_0),
    .Q(main_crg_por_count_TMR_1[5]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52013.11-52019.2" *)
  FD1P3JX \main_crg_por_count_reg[5]_TMR_2  (
    .CK(main_crg_clkout),
    .D(main_crg_por_count_RNO_TMR_2[5]),
    .PD(GND_0),
    .Q(main_crg_por_count_TMR_2[5]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52020.11-52026.2" *)
  FD1P3JX \main_crg_por_count_reg[6]_TMR_0  (
    .CK(main_crg_clkout),
    .D(main_crg_por_count_RNO_TMR_0[6]),
    .PD(GND_0),
    .Q(main_crg_por_count_TMR_0[6]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52020.11-52026.2" *)
  FD1P3JX \main_crg_por_count_reg[6]_TMR_1  (
    .CK(main_crg_clkout),
    .D(main_crg_por_count_RNO_TMR_1[6]),
    .PD(GND_0),
    .Q(main_crg_por_count_TMR_1[6]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52020.11-52026.2" *)
  FD1P3JX \main_crg_por_count_reg[6]_TMR_2  (
    .CK(main_crg_clkout),
    .D(main_crg_por_count_RNO_TMR_2[6]),
    .PD(GND_0),
    .Q(main_crg_por_count_TMR_2[6]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52027.11-52033.2" *)
  FD1P3JX \main_crg_por_count_reg[7]_TMR_0  (
    .CK(main_crg_clkout),
    .D(main_crg_por_count_RNO_TMR_0[7]),
    .PD(GND_0),
    .Q(main_crg_por_count_TMR_0[7]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52027.11-52033.2" *)
  FD1P3JX \main_crg_por_count_reg[7]_TMR_1  (
    .CK(main_crg_clkout),
    .D(main_crg_por_count_RNO_TMR_1[7]),
    .PD(GND_0),
    .Q(main_crg_por_count_TMR_1[7]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52027.11-52033.2" *)
  FD1P3JX \main_crg_por_count_reg[7]_TMR_2  (
    .CK(main_crg_clkout),
    .D(main_crg_por_count_RNO_TMR_2[7]),
    .PD(GND_0),
    .Q(main_crg_por_count_TMR_2[7]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52034.11-52040.2" *)
  FD1P3JX \main_crg_por_count_reg[8]_TMR_0  (
    .CK(main_crg_clkout),
    .D(main_crg_por_count_RNO_TMR_0[8]),
    .PD(GND_0),
    .Q(main_crg_por_count_TMR_0[8]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52034.11-52040.2" *)
  FD1P3JX \main_crg_por_count_reg[8]_TMR_1  (
    .CK(main_crg_clkout),
    .D(main_crg_por_count_RNO_TMR_1[8]),
    .PD(GND_0),
    .Q(main_crg_por_count_TMR_1[8]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52034.11-52040.2" *)
  FD1P3JX \main_crg_por_count_reg[8]_TMR_2  (
    .CK(main_crg_clkout),
    .D(main_crg_por_count_RNO_TMR_2[8]),
    .PD(GND_0),
    .Q(main_crg_por_count_TMR_2[8]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52041.11-52047.2" *)
  FD1P3JX \main_crg_por_count_reg[9]_TMR_0  (
    .CK(main_crg_clkout),
    .D(main_crg_por_count_RNO_TMR_0[9]),
    .PD(GND_0),
    .Q(main_crg_por_count_TMR_0[9]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52041.11-52047.2" *)
  FD1P3JX \main_crg_por_count_reg[9]_TMR_1  (
    .CK(main_crg_clkout),
    .D(main_crg_por_count_RNO_TMR_1[9]),
    .PD(GND_0),
    .Q(main_crg_por_count_TMR_1[9]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:52041.11-52047.2" *)
  FD1P3JX \main_crg_por_count_reg[9]_TMR_2  (
    .CK(main_crg_clkout),
    .D(main_crg_por_count_RNO_TMR_2[9]),
    .PD(GND_0),
    .Q(main_crg_por_count_TMR_2[9]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56014.8-56020.2" *)
  LUT4 main_crg_por_done_11_cZ_TMR_0 (
    .A(main_crg_por_count_TMR_0[7]),
    .B(main_crg_por_count_TMR_0[8]),
    .C(main_crg_por_count_TMR_0[9]),
    .D(main_crg_por_count_TMR_0[10]),
    .Z(main_crg_por_done_11_TMR_0)
  );
  defparam main_crg_por_done_11_cZ_TMR_0.INIT = "0x0001";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56014.8-56020.2" *)
  LUT4 main_crg_por_done_11_cZ_TMR_1 (
    .A(main_crg_por_count_TMR_1[7]),
    .B(main_crg_por_count_TMR_1[8]),
    .C(main_crg_por_count_TMR_1[9]),
    .D(main_crg_por_count_TMR_1[10]),
    .Z(main_crg_por_done_11_TMR_1)
  );
  defparam main_crg_por_done_11_cZ_TMR_1.INIT = "0x0001";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56014.8-56020.2" *)
  LUT4 main_crg_por_done_11_cZ_TMR_2 (
    .A(main_crg_por_count_TMR_2[7]),
    .B(main_crg_por_count_TMR_2[8]),
    .C(main_crg_por_count_TMR_2[9]),
    .D(main_crg_por_count_TMR_2[10]),
    .Z(main_crg_por_done_11_TMR_2)
  );
  defparam main_crg_por_done_11_cZ_TMR_2.INIT = "0x0001";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55915.8-55921.2" *)
  LUT4 main_crg_por_done_12_cZ_TMR_0 (
    .A(main_crg_por_count_TMR_0[0]),
    .B(main_crg_por_count_TMR_0[15]),
    .C(main_crg_por_done_1_TMR_0),
    .D(main_crg_por_done_9_TMR_0),
    .Z(main_crg_por_done_12_TMR_0)
  );
  defparam main_crg_por_done_12_cZ_TMR_0.INIT = "0x1000";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55915.8-55921.2" *)
  LUT4 main_crg_por_done_12_cZ_TMR_1 (
    .A(main_crg_por_count_TMR_1[0]),
    .B(main_crg_por_count_TMR_1[15]),
    .C(main_crg_por_done_1_TMR_1),
    .D(main_crg_por_done_9_TMR_1),
    .Z(main_crg_por_done_12_TMR_1)
  );
  defparam main_crg_por_done_12_cZ_TMR_1.INIT = "0x1000";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55915.8-55921.2" *)
  LUT4 main_crg_por_done_12_cZ_TMR_2 (
    .A(main_crg_por_count_TMR_2[0]),
    .B(main_crg_por_count_TMR_2[15]),
    .C(main_crg_por_done_1_TMR_2),
    .D(main_crg_por_done_9_TMR_2),
    .Z(main_crg_por_done_12_TMR_2)
  );
  defparam main_crg_por_done_12_cZ_TMR_2.INIT = "0x1000";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55924.8-55930.2" *)
  LUT4 main_crg_por_done_13_cZ_TMR_0 (
    .A(main_crg_por_count_TMR_0[13]),
    .B(main_crg_por_count_TMR_0[14]),
    .C(main_crg_por_done_5_TMR_0),
    .D(main_crg_por_done_11_TMR_0),
    .Z(main_crg_por_done_13_TMR_0)
  );
  defparam main_crg_por_done_13_cZ_TMR_0.INIT = "0x1000";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55924.8-55930.2" *)
  LUT4 main_crg_por_done_13_cZ_TMR_1 (
    .A(main_crg_por_count_TMR_1[13]),
    .B(main_crg_por_count_TMR_1[14]),
    .C(main_crg_por_done_5_TMR_1),
    .D(main_crg_por_done_11_TMR_1),
    .Z(main_crg_por_done_13_TMR_1)
  );
  defparam main_crg_por_done_13_cZ_TMR_1.INIT = "0x1000";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55924.8-55930.2" *)
  LUT4 main_crg_por_done_13_cZ_TMR_2 (
    .A(main_crg_por_count_TMR_2[13]),
    .B(main_crg_por_count_TMR_2[14]),
    .C(main_crg_por_done_5_TMR_2),
    .D(main_crg_por_done_11_TMR_2),
    .Z(main_crg_por_done_13_TMR_2)
  );
  defparam main_crg_por_done_13_cZ_TMR_2.INIT = "0x1000";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56237.8-56243.2" *)
  LUT4 main_crg_por_done_1_cZ_TMR_0 (
    .A(main_crg_por_count_TMR_0[5]),
    .B(main_crg_por_count_TMR_0[6]),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_done_1_TMR_0)
  );
  defparam main_crg_por_done_1_cZ_TMR_0.INIT = "0x1111";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56237.8-56243.2" *)
  LUT4 main_crg_por_done_1_cZ_TMR_1 (
    .A(main_crg_por_count_TMR_1[5]),
    .B(main_crg_por_count_TMR_1[6]),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_done_1_TMR_1)
  );
  defparam main_crg_por_done_1_cZ_TMR_1.INIT = "0x1111";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56237.8-56243.2" *)
  LUT4 main_crg_por_done_1_cZ_TMR_2 (
    .A(main_crg_por_count_TMR_2[5]),
    .B(main_crg_por_count_TMR_2[6]),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_done_1_TMR_2)
  );
  defparam main_crg_por_done_1_cZ_TMR_2.INIT = "0x1111";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56246.8-56252.2" *)
  LUT4 main_crg_por_done_5_cZ_TMR_0 (
    .A(main_crg_por_count_TMR_0[11]),
    .B(main_crg_por_count_TMR_0[12]),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_done_5_TMR_0)
  );
  defparam main_crg_por_done_5_cZ_TMR_0.INIT = "0x1111";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56246.8-56252.2" *)
  LUT4 main_crg_por_done_5_cZ_TMR_1 (
    .A(main_crg_por_count_TMR_1[11]),
    .B(main_crg_por_count_TMR_1[12]),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_done_5_TMR_1)
  );
  defparam main_crg_por_done_5_cZ_TMR_1.INIT = "0x1111";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56246.8-56252.2" *)
  LUT4 main_crg_por_done_5_cZ_TMR_2 (
    .A(main_crg_por_count_TMR_2[11]),
    .B(main_crg_por_count_TMR_2[12]),
    .C(GND_0),
    .D(GND_0),
    .Z(main_crg_por_done_5_TMR_2)
  );
  defparam main_crg_por_done_5_cZ_TMR_2.INIT = "0x1111";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56005.8-56011.2" *)
  LUT4 main_crg_por_done_9_cZ_TMR_0 (
    .A(main_crg_por_count_TMR_0[1]),
    .B(main_crg_por_count_TMR_0[2]),
    .C(main_crg_por_count_TMR_0[3]),
    .D(main_crg_por_count_TMR_0[4]),
    .Z(main_crg_por_done_9_TMR_0)
  );
  defparam main_crg_por_done_9_cZ_TMR_0.INIT = "0x0001";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56005.8-56011.2" *)
  LUT4 main_crg_por_done_9_cZ_TMR_1 (
    .A(main_crg_por_count_TMR_1[1]),
    .B(main_crg_por_count_TMR_1[2]),
    .C(main_crg_por_count_TMR_1[3]),
    .D(main_crg_por_count_TMR_1[4]),
    .Z(main_crg_por_done_9_TMR_1)
  );
  defparam main_crg_por_done_9_cZ_TMR_1.INIT = "0x0001";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56005.8-56011.2" *)
  LUT4 main_crg_por_done_9_cZ_TMR_2 (
    .A(main_crg_por_count_TMR_2[1]),
    .B(main_crg_por_count_TMR_2[2]),
    .C(main_crg_por_count_TMR_2[3]),
    .D(main_crg_por_count_TMR_2[4]),
    .Z(main_crg_por_done_9_TMR_2)
  );
  defparam main_crg_por_done_9_cZ_TMR_2.INIT = "0x0001";
  LUT4 main_cs06_0_RED_VOTER (
    .A(main_cs06_TMR_0),
    .B(main_cs06_TMR_1),
    .C(main_cs06_TMR_2),
    .D(1'h0),
    .Z(main_cs06_0_RED_VOTER_wire)
  );
  defparam main_cs06_0_RED_VOTER.INIT = "0xFCC0";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56023.8-56029.2" *)
  LUT4 main_done_11_cZ_TMR_0 (
    .A(main_count_TMR_0[13]),
    .B(main_count_TMR_0[20]),
    .C(main_count_TMR_0[21]),
    .D(main_count_1_TMR_0),
    .Z(main_done_11_TMR_0)
  );
  defparam main_done_11_cZ_TMR_0.INIT = "0x0001";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56023.8-56029.2" *)
  LUT4 main_done_11_cZ_TMR_1 (
    .A(main_count_TMR_1[13]),
    .B(main_count_TMR_1[20]),
    .C(main_count_TMR_1[21]),
    .D(main_count_1_TMR_1),
    .Z(main_done_11_TMR_1)
  );
  defparam main_done_11_cZ_TMR_1.INIT = "0x0001";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56023.8-56029.2" *)
  LUT4 main_done_11_cZ_TMR_2 (
    .A(main_count_TMR_2[13]),
    .B(main_count_TMR_2[20]),
    .C(main_count_TMR_2[21]),
    .D(main_count_1_TMR_2),
    .Z(main_done_11_TMR_2)
  );
  defparam main_done_11_cZ_TMR_2.INIT = "0x0001";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56032.8-56038.2" *)
  LUT4 main_done_12_cZ_TMR_0 (
    .A(main_count_TMR_0[9]),
    .B(main_count_TMR_0[10]),
    .C(main_count_TMR_0[11]),
    .D(main_count_TMR_0[12]),
    .Z(main_done_12_TMR_0)
  );
  defparam main_done_12_cZ_TMR_0.INIT = "0x0001";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56032.8-56038.2" *)
  LUT4 main_done_12_cZ_TMR_1 (
    .A(main_count_TMR_1[9]),
    .B(main_count_TMR_1[10]),
    .C(main_count_TMR_1[11]),
    .D(main_count_TMR_1[12]),
    .Z(main_done_12_TMR_1)
  );
  defparam main_done_12_cZ_TMR_1.INIT = "0x0001";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56032.8-56038.2" *)
  LUT4 main_done_12_cZ_TMR_2 (
    .A(main_count_TMR_2[9]),
    .B(main_count_TMR_2[10]),
    .C(main_count_TMR_2[11]),
    .D(main_count_TMR_2[12]),
    .Z(main_done_12_TMR_2)
  );
  defparam main_done_12_cZ_TMR_2.INIT = "0x0001";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56041.8-56047.2" *)
  LUT4 main_done_13_cZ_TMR_0 (
    .A(main_count_TMR_0[5]),
    .B(main_count_TMR_0[6]),
    .C(main_count_TMR_0[7]),
    .D(main_count_TMR_0[8]),
    .Z(main_done_13_TMR_0)
  );
  defparam main_done_13_cZ_TMR_0.INIT = "0x0001";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56041.8-56047.2" *)
  LUT4 main_done_13_cZ_TMR_1 (
    .A(main_count_TMR_1[5]),
    .B(main_count_TMR_1[6]),
    .C(main_count_TMR_1[7]),
    .D(main_count_TMR_1[8]),
    .Z(main_done_13_TMR_1)
  );
  defparam main_done_13_cZ_TMR_1.INIT = "0x0001";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56041.8-56047.2" *)
  LUT4 main_done_13_cZ_TMR_2 (
    .A(main_count_TMR_2[5]),
    .B(main_count_TMR_2[6]),
    .C(main_count_TMR_2[7]),
    .D(main_count_TMR_2[8]),
    .Z(main_done_13_TMR_2)
  );
  defparam main_done_13_cZ_TMR_2.INIT = "0x0001";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56050.8-56056.2" *)
  LUT4 main_done_15_cZ_TMR_0 (
    .A(main_count_TMR_0[16]),
    .B(main_count_TMR_0[17]),
    .C(main_count_TMR_0[18]),
    .D(main_count_TMR_0[19]),
    .Z(main_done_15_TMR_0)
  );
  defparam main_done_15_cZ_TMR_0.INIT = "0x0001";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56050.8-56056.2" *)
  LUT4 main_done_15_cZ_TMR_1 (
    .A(main_count_TMR_1[16]),
    .B(main_count_TMR_1[17]),
    .C(main_count_TMR_1[18]),
    .D(main_count_TMR_1[19]),
    .Z(main_done_15_TMR_1)
  );
  defparam main_done_15_cZ_TMR_1.INIT = "0x0001";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56050.8-56056.2" *)
  LUT4 main_done_15_cZ_TMR_2 (
    .A(main_count_TMR_2[16]),
    .B(main_count_TMR_2[17]),
    .C(main_count_TMR_2[18]),
    .D(main_count_TMR_2[19]),
    .Z(main_done_15_TMR_2)
  );
  defparam main_done_15_cZ_TMR_2.INIT = "0x0001";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55933.8-55939.2" *)
  LUT4 main_done_16_cZ_TMR_0 (
    .A(main_count_TMR_0[14]),
    .B(main_count_TMR_0[15]),
    .C(main_done_11_TMR_0),
    .D(GND_0),
    .Z(main_done_16_TMR_0)
  );
  defparam main_done_16_cZ_TMR_0.INIT = "0x1010";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55933.8-55939.2" *)
  LUT4 main_done_16_cZ_TMR_1 (
    .A(main_count_TMR_1[14]),
    .B(main_count_TMR_1[15]),
    .C(main_done_11_TMR_1),
    .D(GND_0),
    .Z(main_done_16_TMR_1)
  );
  defparam main_done_16_cZ_TMR_1.INIT = "0x1010";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55933.8-55939.2" *)
  LUT4 main_done_16_cZ_TMR_2 (
    .A(main_count_TMR_2[14]),
    .B(main_count_TMR_2[15]),
    .C(main_done_11_TMR_2),
    .D(GND_0),
    .Z(main_done_16_TMR_2)
  );
  defparam main_done_16_cZ_TMR_2.INIT = "0x1010";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55942.8-55948.2" *)
  LUT4 main_done_18_cZ_TMR_0 (
    .A(main_count_TMR_0[3]),
    .B(main_count_TMR_0[4]),
    .C(main_done_7_TMR_0),
    .D(main_done_15_TMR_0),
    .Z(main_done_18_TMR_0)
  );
  defparam main_done_18_cZ_TMR_0.INIT = "0x1000";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55942.8-55948.2" *)
  LUT4 main_done_18_cZ_TMR_1 (
    .A(main_count_TMR_1[3]),
    .B(main_count_TMR_1[4]),
    .C(main_done_7_TMR_1),
    .D(main_done_15_TMR_1),
    .Z(main_done_18_TMR_1)
  );
  defparam main_done_18_cZ_TMR_1.INIT = "0x1000";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55942.8-55948.2" *)
  LUT4 main_done_18_cZ_TMR_2 (
    .A(main_count_TMR_2[3]),
    .B(main_count_TMR_2[4]),
    .C(main_done_7_TMR_2),
    .D(main_done_15_TMR_2),
    .Z(main_done_18_TMR_2)
  );
  defparam main_done_18_cZ_TMR_2.INIT = "0x1000";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56255.8-56261.2" *)
  LUT4 main_done_7_cZ_TMR_0 (
    .A(main_count_TMR_0[1]),
    .B(main_count_TMR_0[2]),
    .C(GND_0),
    .D(GND_0),
    .Z(main_done_7_TMR_0)
  );
  defparam main_done_7_cZ_TMR_0.INIT = "0x1111";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56255.8-56261.2" *)
  LUT4 main_done_7_cZ_TMR_1 (
    .A(main_count_TMR_1[1]),
    .B(main_count_TMR_1[2]),
    .C(GND_0),
    .D(GND_0),
    .Z(main_done_7_TMR_1)
  );
  defparam main_done_7_cZ_TMR_1.INIT = "0x1111";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56255.8-56261.2" *)
  LUT4 main_done_7_cZ_TMR_2 (
    .A(main_count_TMR_2[1]),
    .B(main_count_TMR_2[2]),
    .C(GND_0),
    .D(GND_0),
    .Z(main_done_7_TMR_2)
  );
  defparam main_done_7_cZ_TMR_2.INIT = "0x1111";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55862.8-55868.2" *)
  LUT4 main_done_cZ_TMR_0 (
    .A(main_done_12_TMR_0),
    .B(main_done_13_TMR_0),
    .C(main_done_16_TMR_0),
    .D(main_done_18_TMR_0),
    .Z(main_done_TMR_0)
  );
  defparam main_done_cZ_TMR_0.INIT = "0x8000";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55862.8-55868.2" *)
  LUT4 main_done_cZ_TMR_1 (
    .A(main_done_12_TMR_1),
    .B(main_done_13_TMR_1),
    .C(main_done_16_TMR_1),
    .D(main_done_18_TMR_1),
    .Z(main_done_TMR_1)
  );
  defparam main_done_cZ_TMR_1.INIT = "0x8000";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55862.8-55868.2" *)
  LUT4 main_done_cZ_TMR_2 (
    .A(main_done_12_TMR_2),
    .B(main_done_13_TMR_2),
    .C(main_done_16_TMR_2),
    .D(main_done_18_TMR_2),
    .Z(main_done_TMR_2)
  );
  defparam main_done_cZ_TMR_2.INIT = "0x8000";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51571.8-51577.2" *)
  LUT4 \main_mode.fb_TMR_0  (
    .A(main_mode_TMR_0),
    .B(main_re_TMR_0),
    .C(GND_0),
    .D(GND_0),
    .Z(\main_mode.fb_0_TMR_0 )
  );
  defparam \main_mode.fb_TMR_0 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51571.8-51577.2" *)
  LUT4 \main_mode.fb_TMR_1  (
    .A(main_mode_TMR_1),
    .B(main_re_TMR_1),
    .C(GND_0),
    .D(GND_0),
    .Z(\main_mode.fb_0_TMR_1 )
  );
  defparam \main_mode.fb_TMR_1 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51571.8-51577.2" *)
  LUT4 \main_mode.fb_TMR_2  (
    .A(main_mode_TMR_2),
    .B(main_re_TMR_2),
    .C(GND_0),
    .D(GND_0),
    .Z(\main_mode.fb_0_TMR_2 )
  );
  defparam \main_mode.fb_TMR_2 .INIT = "0xEEEE";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51971.11-51977.2" *)
  FD1P3IX main_mode_reg_TMR_0 (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(\main_mode.fb_0_TMR_0 ),
    .Q(main_mode_TMR_0),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51971.11-51977.2" *)
  FD1P3IX main_mode_reg_TMR_1 (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(\main_mode.fb_0_TMR_1 ),
    .Q(main_mode_TMR_1),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51971.11-51977.2" *)
  FD1P3IX main_mode_reg_TMR_2 (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(\main_mode.fb_0_TMR_2 ),
    .Q(main_mode_TMR_2),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51964.11-51970.2" *)
  FD1P3IX main_re_reg_TMR_0 (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_storage_0_sqmuxa_TMR_0),
    .Q(main_re_TMR_0),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51964.11-51970.2" *)
  FD1P3IX main_re_reg_TMR_1 (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_storage_0_sqmuxa_TMR_1),
    .Q(main_re_TMR_1),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51964.11-51970.2" *)
  FD1P3IX main_re_reg_TMR_2 (
    .CD(GND_0),
    .CK(sys_clk),
    .D(main_storage_0_sqmuxa_TMR_2),
    .Q(main_re_TMR_2),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51866.11-51872.2" *)
  FD1P3IX \main_storage_reg[0]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[0]),
    .Q(main_storage_TMR_0[0]),
    .SP(builder_csr_bankarray_csrbank1_out0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51866.11-51872.2" *)
  FD1P3IX \main_storage_reg[0]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[0]),
    .Q(main_storage_TMR_1[0]),
    .SP(builder_csr_bankarray_csrbank1_out0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51866.11-51872.2" *)
  FD1P3IX \main_storage_reg[0]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[0]),
    .Q(main_storage_TMR_2[0]),
    .SP(builder_csr_bankarray_csrbank1_out0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51936.11-51942.2" *)
  FD1P3IX \main_storage_reg[10]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[10]),
    .Q(main_storage_TMR_0[10]),
    .SP(builder_csr_bankarray_csrbank1_out0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51936.11-51942.2" *)
  FD1P3IX \main_storage_reg[10]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[10]),
    .Q(main_storage_TMR_1[10]),
    .SP(builder_csr_bankarray_csrbank1_out0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51936.11-51942.2" *)
  FD1P3IX \main_storage_reg[10]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[10]),
    .Q(main_storage_TMR_2[10]),
    .SP(builder_csr_bankarray_csrbank1_out0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51943.11-51949.2" *)
  FD1P3IX \main_storage_reg[11]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[11]),
    .Q(main_storage_TMR_0[11]),
    .SP(builder_csr_bankarray_csrbank1_out0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51943.11-51949.2" *)
  FD1P3IX \main_storage_reg[11]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[11]),
    .Q(main_storage_TMR_1[11]),
    .SP(builder_csr_bankarray_csrbank1_out0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51943.11-51949.2" *)
  FD1P3IX \main_storage_reg[11]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[11]),
    .Q(main_storage_TMR_2[11]),
    .SP(builder_csr_bankarray_csrbank1_out0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51950.11-51956.2" *)
  FD1P3IX \main_storage_reg[12]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[12]),
    .Q(main_storage_TMR_0[12]),
    .SP(builder_csr_bankarray_csrbank1_out0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51950.11-51956.2" *)
  FD1P3IX \main_storage_reg[12]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[12]),
    .Q(main_storage_TMR_1[12]),
    .SP(builder_csr_bankarray_csrbank1_out0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51950.11-51956.2" *)
  FD1P3IX \main_storage_reg[12]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[12]),
    .Q(main_storage_TMR_2[12]),
    .SP(builder_csr_bankarray_csrbank1_out0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51957.11-51963.2" *)
  FD1P3IX \main_storage_reg[13]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[13]),
    .Q(main_storage_TMR_0[13]),
    .SP(builder_csr_bankarray_csrbank1_out0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51957.11-51963.2" *)
  FD1P3IX \main_storage_reg[13]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[13]),
    .Q(main_storage_TMR_1[13]),
    .SP(builder_csr_bankarray_csrbank1_out0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51957.11-51963.2" *)
  FD1P3IX \main_storage_reg[13]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[13]),
    .Q(main_storage_TMR_2[13]),
    .SP(builder_csr_bankarray_csrbank1_out0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51873.11-51879.2" *)
  FD1P3IX \main_storage_reg[1]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[1]),
    .Q(main_storage_TMR_0[1]),
    .SP(builder_csr_bankarray_csrbank1_out0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51873.11-51879.2" *)
  FD1P3IX \main_storage_reg[1]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[1]),
    .Q(main_storage_TMR_1[1]),
    .SP(builder_csr_bankarray_csrbank1_out0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51873.11-51879.2" *)
  FD1P3IX \main_storage_reg[1]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[1]),
    .Q(main_storage_TMR_2[1]),
    .SP(builder_csr_bankarray_csrbank1_out0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51880.11-51886.2" *)
  FD1P3IX \main_storage_reg[2]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[2]),
    .Q(main_storage_TMR_0[2]),
    .SP(builder_csr_bankarray_csrbank1_out0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51880.11-51886.2" *)
  FD1P3IX \main_storage_reg[2]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[2]),
    .Q(main_storage_TMR_1[2]),
    .SP(builder_csr_bankarray_csrbank1_out0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51880.11-51886.2" *)
  FD1P3IX \main_storage_reg[2]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[2]),
    .Q(main_storage_TMR_2[2]),
    .SP(builder_csr_bankarray_csrbank1_out0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51887.11-51893.2" *)
  FD1P3IX \main_storage_reg[3]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[3]),
    .Q(main_storage_TMR_0[3]),
    .SP(builder_csr_bankarray_csrbank1_out0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51887.11-51893.2" *)
  FD1P3IX \main_storage_reg[3]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[3]),
    .Q(main_storage_TMR_1[3]),
    .SP(builder_csr_bankarray_csrbank1_out0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51887.11-51893.2" *)
  FD1P3IX \main_storage_reg[3]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[3]),
    .Q(main_storage_TMR_2[3]),
    .SP(builder_csr_bankarray_csrbank1_out0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51894.11-51900.2" *)
  FD1P3IX \main_storage_reg[4]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[4]),
    .Q(main_storage_TMR_0[4]),
    .SP(builder_csr_bankarray_csrbank1_out0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51894.11-51900.2" *)
  FD1P3IX \main_storage_reg[4]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[4]),
    .Q(main_storage_TMR_1[4]),
    .SP(builder_csr_bankarray_csrbank1_out0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51894.11-51900.2" *)
  FD1P3IX \main_storage_reg[4]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[4]),
    .Q(main_storage_TMR_2[4]),
    .SP(builder_csr_bankarray_csrbank1_out0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51901.11-51907.2" *)
  FD1P3IX \main_storage_reg[5]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[5]),
    .Q(main_storage_TMR_0[5]),
    .SP(builder_csr_bankarray_csrbank1_out0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51901.11-51907.2" *)
  FD1P3IX \main_storage_reg[5]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[5]),
    .Q(main_storage_TMR_1[5]),
    .SP(builder_csr_bankarray_csrbank1_out0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51901.11-51907.2" *)
  FD1P3IX \main_storage_reg[5]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[5]),
    .Q(main_storage_TMR_2[5]),
    .SP(builder_csr_bankarray_csrbank1_out0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51908.11-51914.2" *)
  FD1P3IX \main_storage_reg[6]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[6]),
    .Q(main_storage_TMR_0[6]),
    .SP(builder_csr_bankarray_csrbank1_out0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51908.11-51914.2" *)
  FD1P3IX \main_storage_reg[6]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[6]),
    .Q(main_storage_TMR_1[6]),
    .SP(builder_csr_bankarray_csrbank1_out0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51908.11-51914.2" *)
  FD1P3IX \main_storage_reg[6]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[6]),
    .Q(main_storage_TMR_2[6]),
    .SP(builder_csr_bankarray_csrbank1_out0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51915.11-51921.2" *)
  FD1P3IX \main_storage_reg[7]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[7]),
    .Q(main_storage_TMR_0[7]),
    .SP(builder_csr_bankarray_csrbank1_out0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51915.11-51921.2" *)
  FD1P3IX \main_storage_reg[7]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[7]),
    .Q(main_storage_TMR_1[7]),
    .SP(builder_csr_bankarray_csrbank1_out0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51915.11-51921.2" *)
  FD1P3IX \main_storage_reg[7]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[7]),
    .Q(main_storage_TMR_2[7]),
    .SP(builder_csr_bankarray_csrbank1_out0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51922.11-51928.2" *)
  FD1P3IX \main_storage_reg[8]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[8]),
    .Q(main_storage_TMR_0[8]),
    .SP(builder_csr_bankarray_csrbank1_out0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51922.11-51928.2" *)
  FD1P3IX \main_storage_reg[8]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[8]),
    .Q(main_storage_TMR_1[8]),
    .SP(builder_csr_bankarray_csrbank1_out0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51922.11-51928.2" *)
  FD1P3IX \main_storage_reg[8]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[8]),
    .Q(main_storage_TMR_2[8]),
    .SP(builder_csr_bankarray_csrbank1_out0_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51929.11-51935.2" *)
  FD1P3IX \main_storage_reg[9]_TMR_0  (
    .CD(sys_rst_TMR_0),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_0[9]),
    .Q(main_storage_TMR_0[9]),
    .SP(builder_csr_bankarray_csrbank1_out0_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51929.11-51935.2" *)
  FD1P3IX \main_storage_reg[9]_TMR_1  (
    .CD(sys_rst_TMR_1),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_1[9]),
    .Q(main_storage_TMR_1[9]),
    .SP(builder_csr_bankarray_csrbank1_out0_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51929.11-51935.2" *)
  FD1P3IX \main_storage_reg[9]_TMR_2  (
    .CD(sys_rst_TMR_2),
    .CK(sys_clk),
    .D(dsp_join_kb_0_TMR_2[9]),
    .Q(main_storage_TMR_2[9]),
    .SP(builder_csr_bankarray_csrbank1_out0_re_TMR_2)
  );
  LUT4 main_wren0_0_RED_VOTER (
    .A(main_wren0_TMR_0),
    .B(main_wren0_TMR_1),
    .C(main_wren0_TMR_2),
    .D(1'h0),
    .Z(main_wren0_0_RED_VOTER_wire)
  );
  defparam main_wren0_0_RED_VOTER.INIT = "0xFCC0";
  LUT4 main_wren1_0_RED_VOTER (
    .A(main_wren1_TMR_0),
    .B(main_wren1_TMR_1),
    .C(main_wren1_TMR_2),
    .D(1'h0),
    .Z(main_wren1_0_RED_VOTER_wire)
  );
  defparam main_wren1_0_RED_VOTER.INIT = "0xFCC0";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51819.11-51825.2" *)
  FD1P3IX \mem_adr0_reg[0]_TMR_0  (
    .CD(builder_basesoc_state_TMR_0),
    .CK(sys_clk),
    .D(builder_basesoc_adr_TMR_0[0]),
    .Q(mem_adr0_TMR_0[0]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51819.11-51825.2" *)
  FD1P3IX \mem_adr0_reg[0]_TMR_1  (
    .CD(builder_basesoc_state_TMR_1),
    .CK(sys_clk),
    .D(builder_basesoc_adr_TMR_1[0]),
    .Q(mem_adr0_TMR_1[0]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51819.11-51825.2" *)
  FD1P3IX \mem_adr0_reg[0]_TMR_2  (
    .CD(builder_basesoc_state_TMR_2),
    .CK(sys_clk),
    .D(builder_basesoc_adr_TMR_2[0]),
    .Q(mem_adr0_TMR_2[0]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51827.11-51833.2" *)
  FD1P3IX \mem_adr0_reg[1]_TMR_0  (
    .CD(builder_basesoc_state_TMR_0),
    .CK(sys_clk),
    .D(builder_basesoc_adr_TMR_0[1]),
    .Q(mem_adr0_TMR_0[1]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51827.11-51833.2" *)
  FD1P3IX \mem_adr0_reg[1]_TMR_1  (
    .CD(builder_basesoc_state_TMR_1),
    .CK(sys_clk),
    .D(builder_basesoc_adr_TMR_1[1]),
    .Q(mem_adr0_TMR_1[1]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51827.11-51833.2" *)
  FD1P3IX \mem_adr0_reg[1]_TMR_2  (
    .CD(builder_basesoc_state_TMR_2),
    .CK(sys_clk),
    .D(builder_basesoc_adr_TMR_2[1]),
    .Q(mem_adr0_TMR_2[1]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51835.11-51841.2" *)
  FD1P3IX \mem_adr0_reg[2]_TMR_0  (
    .CD(builder_basesoc_state_TMR_0),
    .CK(sys_clk),
    .D(builder_basesoc_adr_TMR_0[2]),
    .Q(mem_adr0_TMR_0[2]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51835.11-51841.2" *)
  FD1P3IX \mem_adr0_reg[2]_TMR_1  (
    .CD(builder_basesoc_state_TMR_1),
    .CK(sys_clk),
    .D(builder_basesoc_adr_TMR_1[2]),
    .Q(mem_adr0_TMR_1[2]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51835.11-51841.2" *)
  FD1P3IX \mem_adr0_reg[2]_TMR_2  (
    .CD(builder_basesoc_state_TMR_2),
    .CK(sys_clk),
    .D(builder_basesoc_adr_TMR_2[2]),
    .Q(mem_adr0_TMR_2[2]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51843.11-51849.2" *)
  FD1P3IX \mem_adr0_reg[3]_TMR_0  (
    .CD(builder_basesoc_state_TMR_0),
    .CK(sys_clk),
    .D(builder_basesoc_adr_TMR_0[3]),
    .Q(mem_adr0_TMR_0[3]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51843.11-51849.2" *)
  FD1P3IX \mem_adr0_reg[3]_TMR_1  (
    .CD(builder_basesoc_state_TMR_1),
    .CK(sys_clk),
    .D(builder_basesoc_adr_TMR_1[3]),
    .Q(mem_adr0_TMR_1[3]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51843.11-51849.2" *)
  FD1P3IX \mem_adr0_reg[3]_TMR_2  (
    .CD(builder_basesoc_state_TMR_2),
    .CK(sys_clk),
    .D(builder_basesoc_adr_TMR_2[3]),
    .Q(mem_adr0_TMR_2[3]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51851.11-51857.2" *)
  FD1P3IX \mem_adr0_reg[4]_TMR_0  (
    .CD(builder_basesoc_state_TMR_0),
    .CK(sys_clk),
    .D(builder_basesoc_adr_TMR_0[4]),
    .Q(mem_adr0_TMR_0[4]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51851.11-51857.2" *)
  FD1P3IX \mem_adr0_reg[4]_TMR_1  (
    .CD(builder_basesoc_state_TMR_1),
    .CK(sys_clk),
    .D(builder_basesoc_adr_TMR_1[4]),
    .Q(mem_adr0_TMR_1[4]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51851.11-51857.2" *)
  FD1P3IX \mem_adr0_reg[4]_TMR_2  (
    .CD(builder_basesoc_state_TMR_2),
    .CK(sys_clk),
    .D(builder_basesoc_adr_TMR_2[4]),
    .Q(mem_adr0_TMR_2[4]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51859.11-51865.2" *)
  FD1P3IX \mem_adr0_reg[5]_TMR_0  (
    .CD(builder_basesoc_state_TMR_0),
    .CK(sys_clk),
    .D(builder_basesoc_adr_TMR_0[5]),
    .Q(mem_adr0_TMR_0[5]),
    .SP(VCC_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51859.11-51865.2" *)
  FD1P3IX \mem_adr0_reg[5]_TMR_1  (
    .CD(builder_basesoc_state_TMR_1),
    .CK(sys_clk),
    .D(builder_basesoc_adr_TMR_1[5]),
    .Q(mem_adr0_TMR_1[5]),
    .SP(VCC_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51859.11-51865.2" *)
  FD1P3IX \mem_adr0_reg[5]_TMR_2  (
    .CD(builder_basesoc_state_TMR_2),
    .CK(sys_clk),
    .D(builder_basesoc_adr_TMR_2[5]),
    .Q(mem_adr0_TMR_2[5]),
    .SP(VCC_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:59198.9-59207.2" *)
  SP16K rom_dat0_2_0_0 (
    .AD({ builder_array_muxed0_12_RED_VOTER_wire, builder_array_muxed0_11_RED_VOTER_wire, builder_array_muxed0_10_RED_VOTER_wire, builder_array_muxed0_9_RED_VOTER_wire, builder_array_muxed0_8_RED_VOTER_wire, builder_array_muxed0_7_RED_VOTER_wire, builder_array_muxed0_6_RED_VOTER_wire, builder_array_muxed0_5_RED_VOTER_wire, builder_array_muxed0_4_RED_VOTER_wire, N_103_0_RED_VOTER_wire, builder_array_muxed0_2_RED_VOTER_wire, builder_array_muxed0_1_RED_VOTER_wire, builder_array_muxed0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire }),
    .CE(VCC_0_RED_VOTER_wire),
    .CLK(sys_clk),
    .CS({ VCC_0_RED_VOTER_wire, VCC_0_RED_VOTER_wire, VCC_0_RED_VOTER_wire }),
    .DI({ GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire }),
    .DO({ rom_dat0_2_0_0_DO, rom_dat0[1:0] }),
    .RST(GND_0_0_RED_VOTER_wire),
    .WE(GND_0_0_RED_VOTER_wire)
  );
  defparam rom_dat0_2_0_0.DATA_WIDTH = "X2";
  defparam rom_dat0_2_0_0.GSR = "ENABLED";
  defparam rom_dat0_2_0_0.INITVAL_00 = "0x3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF";
  defparam rom_dat0_2_0_0.INITVAL_01 = "0x3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF";
  defparam rom_dat0_2_0_0.INITVAL_02 = "0x3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF";
  defparam rom_dat0_2_0_0.INITVAL_03 = "0x3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF";
  defparam rom_dat0_2_0_0.INITVAL_04 = "0x3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF";
  defparam rom_dat0_2_0_0.INITVAL_05 = "0x3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF";
  defparam rom_dat0_2_0_0.INITVAL_06 = "0x3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF";
  defparam rom_dat0_2_0_0.INITVAL_07 = "0x3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF";
  defparam rom_dat0_2_0_0.INITVAL_08 = "0x3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF";
  defparam rom_dat0_2_0_0.INITVAL_09 = "0x3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF";
  defparam rom_dat0_2_0_0.INITVAL_0A = "0x3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF";
  defparam rom_dat0_2_0_0.INITVAL_0B = "0x3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF";
  defparam rom_dat0_2_0_0.INITVAL_0C = "0x3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF";
  defparam rom_dat0_2_0_0.INITVAL_0D = "0x3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF";
  defparam rom_dat0_2_0_0.INITVAL_0E = "0x3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF";
  defparam rom_dat0_2_0_0.INITVAL_0F = "0x3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF";
  defparam rom_dat0_2_0_0.INITVAL_10 = "0x3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF";
  defparam rom_dat0_2_0_0.INITVAL_11 = "0x3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF";
  defparam rom_dat0_2_0_0.INITVAL_12 = "0x3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF";
  defparam rom_dat0_2_0_0.INITVAL_13 = "0x3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF";
  defparam rom_dat0_2_0_0.INITVAL_14 = "0x3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF";
  defparam rom_dat0_2_0_0.INITVAL_15 = "0x3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF";
  defparam rom_dat0_2_0_0.INITVAL_16 = "0x3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF";
  defparam rom_dat0_2_0_0.INITVAL_17 = "0x3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF";
  defparam rom_dat0_2_0_0.INITVAL_18 = "0x3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF";
  defparam rom_dat0_2_0_0.INITVAL_19 = "0x3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF";
  defparam rom_dat0_2_0_0.INITVAL_1A = "0x3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF";
  defparam rom_dat0_2_0_0.INITVAL_1B = "0x3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF";
  defparam rom_dat0_2_0_0.INITVAL_1C = "0x3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF";
  defparam rom_dat0_2_0_0.INITVAL_1D = "0x3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF";
  defparam rom_dat0_2_0_0.INITVAL_1E = "0x3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF";
  defparam rom_dat0_2_0_0.INITVAL_1F = "0x3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF";
  defparam rom_dat0_2_0_0.INITVAL_20 = "0x3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF";
  defparam rom_dat0_2_0_0.INITVAL_21 = "0x1240B3FC24264543CC55200CF14CFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF3FCFF";
  defparam rom_dat0_2_0_0.INITVAL_22 = "0x1205210C023209C0906830C1C0900305C6B044641C05030000104F003CC601021270EF0C4CC38C0C";
  defparam rom_dat0_2_0_0.INITVAL_23 = "0x2002011009024882342109C270904C0D825094ED0C4D0020C0010000A4141500036411030342DCC4";
  defparam rom_dat0_2_0_0.INITVAL_24 = "0x040070882531C7708C371C0043C036394F508844124501E00D130041F80C090760EC6D0EC4020000";
  defparam rom_dat0_2_0_0.INITVAL_25 = "0x104421B4DC0480405C20100C6284333FC0C0F0C32CCC00EC0C30C1422CB8090B7024090244E308F5";
  defparam rom_dat0_2_0_0.INITVAL_26 = "0x0000F3FCFF3FCFF04412278B73545F3D45B1785514415188FC378D11FC32078CB204FC1945535457";
  defparam rom_dat0_2_0_0.INITVAL_27 = "0x0180030000000000000000000008AA204551000000000000C4130441208801048220000000000000";
  defparam rom_dat0_2_0_0.INITVAL_28 = "0x34C9324C932B06C1B06C1E4390E439018C6318C634C9324C932B06C1B06C1E4390E4390000000000";
  defparam rom_dat0_2_0_0.INITVAL_29 = "0x34C9324C932B06C1B06C1E4390E439018C6318C634C9324C932B06C1B06C1E4390E439018C6318C6";
  defparam rom_dat0_2_0_0.INITVAL_2A = "0x074C82DC62074C82DC62074C82DC62074C82DC62074C82DC62074C82DC62074C82DC62018C6318C6";
  defparam rom_dat0_2_0_0.INITVAL_2B = "0x074C82DC62074C82DC62074C82DC62074C82DC62074C82DC62074C82DC62074C82DC62074C82DC62";
  defparam rom_dat0_2_0_0.INITVAL_2C = "0x00000000000000000C5D10C800E0022C05434C34244732101101036008D50001515454174C82DC62";
  defparam rom_dat0_2_0_0.INITVAL_2D = "0x37CF0000000000000C0000C0000C0000C0000C0000C0000C40100402008020080200802000000000";
  defparam rom_dat0_2_0_0.INITVAL_2E = "0x0000000000000000000000000000000000000000000000000000000000000000000C000000030000";
  defparam rom_dat0_2_0_0.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_0.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_0.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_0.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_0.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_0.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_0.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_0.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_0.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_0.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_0.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_0.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_0.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_0.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_0.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_0.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_0.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_0.OUTREG = "BYPASSED";
  defparam rom_dat0_2_0_0.RESETMODE = "SYNC";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:59117.9-59126.2" *)
  SP16K rom_dat0_2_0_1 (
    .AD({ builder_array_muxed0_12_RED_VOTER_wire, builder_array_muxed0_11_RED_VOTER_wire, builder_array_muxed0_10_RED_VOTER_wire, builder_array_muxed0_9_RED_VOTER_wire, builder_array_muxed0_8_RED_VOTER_wire, builder_array_muxed0_7_RED_VOTER_wire, builder_array_muxed0_6_RED_VOTER_wire, builder_array_muxed0_5_RED_VOTER_wire, builder_array_muxed0_4_RED_VOTER_wire, N_103_0_RED_VOTER_wire, builder_array_muxed0_2_RED_VOTER_wire, builder_array_muxed0_1_RED_VOTER_wire, builder_array_muxed0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire }),
    .CE(VCC_0_RED_VOTER_wire),
    .CLK(sys_clk),
    .CS({ VCC_0_RED_VOTER_wire, VCC_0_RED_VOTER_wire, VCC_0_RED_VOTER_wire }),
    .DI({ GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire }),
    .DO({ rom_dat0_2_0_1_DO, rom_dat0[3:2] }),
    .RST(GND_0_0_RED_VOTER_wire),
    .WE(GND_0_0_RED_VOTER_wire)
  );
  defparam rom_dat0_2_0_1.DATA_WIDTH = "X2";
  defparam rom_dat0_2_0_1.GSR = "ENABLED";
  defparam rom_dat0_2_0_1.INITVAL_00 = "0x1000000000000000000000000000011401F01C0011C000104404400000000000C000000000000003";
  defparam rom_dat0_2_0_1.INITVAL_01 = "0x000000C0003000004000300C300000000000C000000000000000C00000000C000030003000000000";
  defparam rom_dat0_2_0_1.INITVAL_02 = "0x00C0000003030C0000000000000C000000000000000C030000300000000000003000000003000000";
  defparam rom_dat0_2_0_1.INITVAL_03 = "0x0C03C0000C0000C00041000030F0F100004000041001C1C0000001F000F000C0331C0000401000C0";
  defparam rom_dat0_2_0_1.INITVAL_04 = "0x014740000001000130C730C00000000CCCC0000000010000000C0030FC100C0C0000000000C0CCCC";
  defparam rom_dat0_2_0_1.INITVAL_05 = "0x000400000000C310000000C040C04C0400C00004330F30CC00000C00003000C00130100301000000";
  defparam rom_dat0_2_0_1.INITVAL_06 = "0x1100000001040000000C000C00003011070000140107D010000044031000004000C0300000005007";
  defparam rom_dat0_2_0_1.INITVAL_07 = "0x030040000C100300000003043010C01F04C31003004003100300000310313104031003000030440C";
  defparam rom_dat0_2_0_1.INITVAL_08 = "0x00000310300000C10030000C400C010000C10030000000C40C1C0C303000000003000C1003000C10";
  defparam rom_dat0_2_0_1.INITVAL_09 = "0x00C000000C13C030400C00040030400C000000C431C4304000300030400C030400C01000031000C0";
  defparam rom_dat0_2_0_1.INITVAL_0A = "0x000C000000310413C00C1003000C10030000C40030040000C400C00000003103C0C40030004000C4";
  defparam rom_dat0_2_0_1.INITVAL_0B = "0x01C070005C014C70C4CF070C7070C70707131C34000003000C10030000C400C000C4003000400031";
  defparam rom_dat0_2_0_1.INITVAL_0C = "0x000000C03001000000000000007000140000000000010040F030C0300C0301C053C4CC13C1F0CC07";
  defparam rom_dat0_2_0_1.INITVAL_0D = "0x000010000000000300000000000000030F007C000C0000100C000000003000C1000400000C00C033";
  defparam rom_dat0_2_0_1.INITVAL_0E = "0x0000000030000001C0C000C00000000001005000110410700C0001330400000040300004C0000003";
  defparam rom_dat0_2_0_1.INITVAL_0F = "0x0C00C014F000000000300000300C0C0C013000C0000003C000000400000300C00300001040010000";
  defparam rom_dat0_2_0_1.INITVAL_10 = "0x0000030C3304003300F00C0000000300C030003004C000000C0C00C0300004000000030003030030";
  defparam rom_dat0_2_0_1.INITVAL_11 = "0x000010F00C0303000C300000C0000000040000410F000040400001C300C00C013000003C00003000";
  defparam rom_dat0_2_0_1.INITVAL_12 = "0x010010CC0300C000C000000000000000000000000000010440000040000000C1C310010004003001";
  defparam rom_dat0_2_0_1.INITVAL_13 = "0x0000030400010010004C00000010400000000C10000C100000010C100000010410040305C0300400";
  defparam rom_dat0_2_0_1.INITVAL_14 = "0x0000000000000000C00300000000000000000C100000410000000000503000000040C10100000000";
  defparam rom_dat0_2_0_1.INITVAL_15 = "0x0C00300030030300000C0300000C3303001000000000000000304000000000001044000000000004";
  defparam rom_dat0_2_0_1.INITVAL_16 = "0x0300C0C00000000000000000004000000000040030000040C30000000C0000C3000000000000000C";
  defparam rom_dat0_2_0_1.INITVAL_17 = "0x00C030C0430001D000C0100300000000010000000000000000004000000000000000000000C0C000";
  defparam rom_dat0_2_0_1.INITVAL_18 = "0x030C100004000100001000000000400003004031000C40300000031000030C0040C0CC00C0C30C00";
  defparam rom_dat0_2_0_1.INITVAL_19 = "0x00003030400000000030000000C00000C0000C0C3300000C00000300300000000000001003003001";
  defparam rom_dat0_2_0_1.INITVAL_1A = "0x000000000400000000000000000040004C00C000000C30C00000C000000000000000000000000000";
  defparam rom_dat0_2_0_1.INITVAL_1B = "0x000000000000000000000000000000004000000004000000001C00000010004100300C1000000000";
  defparam rom_dat0_2_0_1.INITVAL_1C = "0x04000040011C0430C04000C10000C4000070400131004100040C4000001031000000411C00000000";
  defparam rom_dat0_2_0_1.INITVAL_1D = "0x3300000001000000000000000014F00000004070000C00C00030010000133001001CC00001104030";
  defparam rom_dat0_2_0_1.INITVAL_1E = "0x100000303000010000000C0CC0000300C100000000031300410003731C040401000000000000004C";
  defparam rom_dat0_2_0_1.INITVAL_1F = "0x0004000C0003000330701000031CC0004C0110000007F0707C0001C010400000000007070C430000";
  defparam rom_dat0_2_0_1.INITVAL_20 = "0x04C0000040014440700000000054140007305000000313007007004000C0030030101000033070C0";
  defparam rom_dat0_2_0_1.INITVAL_21 = "0x364033303818CFC2F8FF2804D144C00101110000110441C40C000410000010005000540300004010";
  defparam rom_dat0_2_0_1.INITVAL_22 = "0x1901913030034211287308023120CC1906F3886C3D854140801080020007010210F46E1140D10C10";
  defparam rom_dat0_2_0_1.INITVAL_23 = "0x3C06435452148F30CC01120701204103849124B9314700100800000028370640805466004B001001";
  defparam rom_dat0_2_0_1.INITVAL_24 = "0x38C3C0000C0545C0000C0C41D0C44F3300D0D083048C30A0531A41E1387103045310FF310E93C069";
  defparam rom_dat0_2_0_1.INITVAL_25 = "0x22842114E00002802C02200B4004233FC080F0C22BCE00A80C3083C00C330303004812048C804019";
  defparam rom_dat0_2_0_1.INITVAL_26 = "0x364AA2A8AA2BCFF04415308EA2FCFB0BCFB1FCFF3DC3F398882A083288100A0812488827CFF03CFD";
  defparam rom_dat0_2_0_1.INITVAL_27 = "0x2C8E80000000000000000000000000000000044000008024472B4070844F094031B40C0000B20418";
  defparam rom_dat0_2_0_1.INITVAL_28 = "0x1A8BF300151A8BF300151A8BF300151FCEA254400FCEA254400FCEA254400FCEA254400686A2A8AE";
  defparam rom_dat0_2_0_1.INITVAL_29 = "0x300151A8BF300151A8BF300151A8BF354400FCEA254400FCEA254400FCEA254400FCEA2A8BF30015";
  defparam rom_dat0_2_0_1.INITVAL_2A = "0x3B4072B407248F8148F811CAD01CAD0E0523E0523B4072B407248F8148F811CAD01CAD000151A8BF";
  defparam rom_dat0_2_0_1.INITVAL_2B = "0x3B4072B407248F8148F811CAD01CAD0E0523E0523B4072B407248F8148F811CAD01CAD0E0523E052";
  defparam rom_dat0_2_0_1.INITVAL_2C = "0x0480900000000033CC7935011104160001D04C482804301031020072000700099194941E0523E052";
  defparam rom_dat0_2_0_1.INITVAL_2D = "0x03CF00000021400000000000000000000000000000000000340D03201C0401406018070DC3408C0F";
  defparam rom_dat0_2_0_1.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000008050000000000";
  defparam rom_dat0_2_0_1.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_1.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_1.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_1.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_1.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_1.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_1.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_1.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_1.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_1.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_1.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_1.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_1.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_1.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_1.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_1.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_1.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_1.OUTREG = "BYPASSED";
  defparam rom_dat0_2_0_1.RESETMODE = "SYNC";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:58388.9-58397.2" *)
  SP16K rom_dat0_2_0_10 (
    .AD({ builder_array_muxed0_12_RED_VOTER_wire, builder_array_muxed0_11_RED_VOTER_wire, builder_array_muxed0_10_RED_VOTER_wire, builder_array_muxed0_9_RED_VOTER_wire, builder_array_muxed0_8_RED_VOTER_wire, builder_array_muxed0_7_RED_VOTER_wire, builder_array_muxed0_6_RED_VOTER_wire, builder_array_muxed0_5_RED_VOTER_wire, builder_array_muxed0_4_RED_VOTER_wire, N_103_0_RED_VOTER_wire, builder_array_muxed0_2_RED_VOTER_wire, builder_array_muxed0_1_RED_VOTER_wire, builder_array_muxed0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire }),
    .CE(VCC_0_RED_VOTER_wire),
    .CLK(sys_clk),
    .CS({ VCC_0_RED_VOTER_wire, VCC_0_RED_VOTER_wire, VCC_0_RED_VOTER_wire }),
    .DI({ GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire }),
    .DO({ rom_dat0_2_0_10_DO, rom_dat0[21:20] }),
    .RST(GND_0_0_RED_VOTER_wire),
    .WE(GND_0_0_RED_VOTER_wire)
  );
  defparam rom_dat0_2_0_10.DATA_WIDTH = "X2";
  defparam rom_dat0_2_0_10.GSR = "ENABLED";
  defparam rom_dat0_2_0_10.INITVAL_00 = "0x0000000003330000345916C9338844000000040C00404300010008000000000003904E138E500000";
  defparam rom_dat0_2_0_10.INITVAL_01 = "0x024C017083140003342910C4D100300D03304029390082F0060148C03C041084D0C060110153F425";
  defparam rom_dat0_2_0_10.INITVAL_02 = "0x0C403070611D84C15C40004702C43C30C003C0C01C04C1703111CF300000220D114CD4144D50005C";
  defparam rom_dat0_2_0_10.INITVAL_03 = "0x3649500C6730007210101600D05440018D029804000000384D210010000000001000440100030C4F";
  defparam rom_dat0_2_0_10.INITVAL_04 = "0x040101043930081010411544903401074760280E00400000001709D2440C1704C308160E00436466";
  defparam rom_dat0_2_0_10.INITVAL_05 = "0x004020E84810054020280040004004000250C00015051144010044F0081100440010010100000000";
  defparam rom_dat0_2_0_10.INITVAL_06 = "0x00031000400000000C54084400100000010190403800400001010101000000000000010001320401";
  defparam rom_dat0_2_0_10.INITVAL_07 = "0x0000000004000021000C110250005005000100000000010000140001085010000100001000102004";
  defparam rom_dat0_2_0_10.INITVAL_08 = "0x10008008950D484000000D8400000000000000093001000094048690546B0108000084000000E400";
  defparam rom_dat0_2_0_10.INITVAL_09 = "0x0006001000090010000003400000000180010002104050080400081000000100000000000000000D";
  defparam rom_dat0_2_0_10.INITVAL_0A = "0x00027000400082414004008000F4002000C24000000000000000027000400085434000000D000000";
  defparam rom_dat0_2_0_10.INITVAL_0B = "0x00000000000C0000000000000000000000000010038441000400010070400040324000100D000000";
  defparam rom_dat0_2_0_10.INITVAL_0C = "0x208000401C000000000003003010E0030000384E120C101050100000040000400040000100000000";
  defparam rom_dat0_2_0_10.INITVAL_0D = "0x0C0000300001C90158C40000023808010500140304004088471042430800004000C0710000414051";
  defparam rom_dat0_2_0_10.INITVAL_0E = "0x378F61B411200F9048633F43400C950C0C8008000080C01C4403C411000000CC31100F000BD0D005";
  defparam rom_dat0_2_0_10.INITVAL_0F = "0x03004000540000401C1030C000C404040013002C3B00F140003340037C753141C00800040020FC13";
  defparam rom_dat0_2_0_10.INITVAL_10 = "0x0003C0045003CC10C04407433030C0310C033000000B12BC070000710038000000003103C001E004";
  defparam rom_dat0_2_0_10.INITVAL_11 = "0x0900804C073001F2841038C0103000048103D03004C340100D310040C030000C12C490130130040C";
  defparam rom_dat0_2_0_10.INITVAL_12 = "0x200D80745D17484374A71B0040500E05C04108450084100022020002202000404180D02803D110E0";
  defparam rom_dat0_2_0_10.INITVAL_13 = "0x2E4181C0C40000C328373402C3000030040064480CC4400C9400044110283001C3A0F10049100070";
  defparam rom_dat0_2_0_10.INITVAL_14 = "0x000000007407800040310007F0C0010D0632440804C030000C208500000109400330700000001000";
  defparam rom_dat0_2_0_10.INITVAL_15 = "0x04009000D00D090000260584230411080440E0B00E892200C010007274430003030022390E724400";
  defparam rom_dat0_2_0_10.INITVAL_16 = "0x01C0104883000322E0003001500000000000C0400802B0004100C0007431074080300D16CC00C094";
  defparam rom_dat0_2_0_10.INITVAL_17 = "0x00401060110080421048044CC00C3F1100000420100383400203080200043000400C0020C5404000";
  defparam rom_dat0_2_0_10.INITVAL_18 = "0x000103840025004150011F0AF340053C01F0101000C4101443020900009D060400486504406104C0";
  defparam rom_dat0_2_0_10.INITVAL_19 = "0x0E01800000000020B8031380300044014102A000180EC074F1010002003000000150E00001438040";
  defparam rom_dat0_2_0_10.INITVAL_1A = "0x29C6D344013A856164390A41C3703807C73040301B80004C171045005C3339C4E34C253EC570C088";
  defparam rom_dat0_2_0_10.INITVAL_1B = "0x3883B2043B0803B20C3B0B00B3700B300FC0ACD030C47020FC074032000E0C000014040989C1985D";
  defparam rom_dat0_2_0_10.INITVAL_1C = "0x00433170C824001050000040022840228C102CBD100B10B8D90500A2500B1402A140200600B2CC0B";
  defparam rom_dat0_2_0_10.INITVAL_1D = "0x1548801C500000524C830D431000400601900C152185925486164800041108412024082142000414";
  defparam rom_dat0_2_0_10.INITVAL_1E = "0x030103105000400000780405401801004400000000010120003041010400230400200E134E604005";
  defparam rom_dat0_2_0_10.INITVAL_1F = "0x3900010400010E411010000001042408C42040080A4110101211834084322A0C826C010104011480";
  defparam rom_dat0_2_0_10.INITVAL_20 = "0x004F43300300002114AC0F4020000012014000000000000800200210204401001000000001101064";
  defparam rom_dat0_2_0_10.INITVAL_21 = "0x28CAB2A48A2A0FF3ACFF0ECBA2804600C00010B800000060C0380002083000C402C00300C3703000";
  defparam rom_dat0_2_0_10.INITVAL_22 = "0x230AB0AC2E038A22A0BE23CAE3A0B8288CE2B4A02B8AA2B83B2A8802AC00230B3280820C88E0ACFA";
  defparam rom_dat0_2_0_10.INITVAL_23 = "0x2ACEA3A8EA3A8EE3B83A3A0AA2A0EA2E0EB2A09B2FCA33FC6E3E4FF308BA2EC882F8A20ACAE2288A";
  defparam rom_dat0_2_0_10.INITVAL_24 = "0x2BC383E82A3A8283EC382EC382EC283A8B82B88E2E86F2FCFA1ACB82B86A2A0EE2ACAE3AC8E2ACEE";
  defparam rom_dat0_2_0_10.INITVAL_25 = "0x3F8A33B8B80ECEA228BE2A0AE3A8B12586C1E86B0DC6A2CC6A2AC332208819C8B0E83A0E83D2A82E";
  defparam rom_dat0_2_0_10.INITVAL_26 = "0x0000F3FC0000000088233AC3A33CFA2FCF22B83F3D87F320CC0A0CA29C0B2A4C10289C2CCFF15CFC";
  defparam rom_dat0_2_0_10.INITVAL_27 = "0x0283100000000000000000000010000100001005168AA28000000000000000000000000000000000";
  defparam rom_dat0_2_0_10.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_10.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_10.INITVAL_2A = "0x0002A2547F3547F3002A2A8800FCD51A8800FCD51547F3002A2002A2547F3FCD51A8800000000000";
  defparam rom_dat0_2_0_10.INITVAL_2B = "0x3FCD51A8800A8800FCD51547F3002A2547F3002A2A8800FCD51FCD51A8800002A2547F3FCD51A880";
  defparam rom_dat0_2_0_10.INITVAL_2C = "0x000000000000000000E3228A82A88A3A8BA2A0A9088F222CA22242E3A8AE088E333C3C3002A2547F";
  defparam rom_dat0_2_0_10.INITVAL_2D = "0x00CF0000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_10.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_10.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_10.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_10.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_10.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_10.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_10.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_10.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_10.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_10.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_10.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_10.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_10.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_10.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_10.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_10.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_10.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_10.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_10.OUTREG = "BYPASSED";
  defparam rom_dat0_2_0_10.RESETMODE = "SYNC";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:58307.9-58316.2" *)
  SP16K rom_dat0_2_0_11 (
    .AD({ builder_array_muxed0_12_RED_VOTER_wire, builder_array_muxed0_11_RED_VOTER_wire, builder_array_muxed0_10_RED_VOTER_wire, builder_array_muxed0_9_RED_VOTER_wire, builder_array_muxed0_8_RED_VOTER_wire, builder_array_muxed0_7_RED_VOTER_wire, builder_array_muxed0_6_RED_VOTER_wire, builder_array_muxed0_5_RED_VOTER_wire, builder_array_muxed0_4_RED_VOTER_wire, N_103_0_RED_VOTER_wire, builder_array_muxed0_2_RED_VOTER_wire, builder_array_muxed0_1_RED_VOTER_wire, builder_array_muxed0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire }),
    .CE(VCC_0_RED_VOTER_wire),
    .CLK(sys_clk),
    .CS({ VCC_0_RED_VOTER_wire, VCC_0_RED_VOTER_wire, VCC_0_RED_VOTER_wire }),
    .DI({ GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire }),
    .DO({ rom_dat0_2_0_11_DO, rom_dat0[23:22] }),
    .RST(GND_0_0_RED_VOTER_wire),
    .WE(GND_0_0_RED_VOTER_wire)
  );
  defparam rom_dat0_2_0_11.DATA_WIDTH = "X2";
  defparam rom_dat0_2_0_11.GSR = "ENABLED";
  defparam rom_dat0_2_0_11.INITVAL_00 = "0x004B12C4B3374003048C0E8A90245A10400104490CC5C2C431200012C4B12C4B43FC0F3E85400000";
  defparam rom_dat0_2_0_11.INITVAL_01 = "0x0C004030D03C03C324C01CC4C0EC71048191A0C020CD00D873108CC37C43340B8398EF300101D0C3";
  defparam rom_dat0_2_0_11.INITVAL_02 = "0x2D431114342F07C00C03330303483617C013D0C10E04D2303C00CFB00CC7020C400800030603100E";
  defparam rom_dat0_2_0_11.INITVAL_03 = "0x01041000200400400C0112091000A000C803CC000088F09452084020380000000100F00A02030C8F";
  defparam rom_dat0_2_0_11.INITVAL_04 = "0x28020260950800203070214E300C200E8AA208720B00306C1B0E05F2E08C0C80C3AC8F2283216421";
  defparam rom_dat0_2_0_11.INITVAL_05 = "0x000030E00C00C200302D000032900C238280C020134640B8AA0104F01C260101103802030C6318C7";
  defparam rom_dat0_2_0_11.INITVAL_06 = "0x0403C100000006C1BC8F010701AC0404002054820000C1006E00028140B12C000050020400400880";
  defparam rom_dat0_2_0_11.INITVAL_07 = "0x0DC102C4BD000C40B0002382208C4C0BC080800E0D01B1400E0B0081C8281400B1400E0B0001203E";
  defparam rom_dat0_2_0_11.INITVAL_08 = "0x0B0001081C0FC01000CC2C090038C40C4BD000C00C02209081090411100A344003CCD1000CC2C440";
  defparam rom_dat0_2_0_11.INITVAL_09 = "0x0380C0208D0980500034370012F400300C0220523C00230050100C2100370900033042318E000CD2";
  defparam rom_dat0_2_0_11.INITVAL_0A = "0x00CC030088108301000B008CC3CC002DC2C050033C40B06C5003840300881082035003334C006C50";
  defparam rom_dat0_2_0_11.INITVAL_0B = "0x300003040D280503A07C03C7013C6013028100D0000A020004000C3380C00383B000033C4C0318E4";
  defparam rom_dat0_2_0_11.INITVAL_0C = "0x24400000C9000C6318C630003010610003C028A40D40D220E3148310C0C2000303A07C010CC3B040";
  defparam rom_dat0_2_0_11.INITVAL_0D = "0x04C1C2B800000280300C0C0030340802028000C80902008C0B0040000840000C10C000000CC0E016";
  defparam rom_dat0_2_0_11.INITVAL_0E = "0x3F8F50B8B5310FA0D8873B47000458120C020C0300C0C01C0F00C001B0312CCC303C03000AC28020";
  defparam rom_dat0_2_0_11.INITVAL_0F = "0x2700E300603000902CE03CC120C0AC28C0C320682B03F08C001380A37CFA18C6008088080380DC3B";
  defparam rom_dat0_2_0_11.INITVAL_10 = "0x000FF1BC2003C8F1E8E0274F3030CD310E833023030A02BC3F3A03B0F03C300312D8F30FCEB0FC22";
  defparam rom_dat0_2_0_11.INITVAL_11 = "0x0C0000FCAB3F8CA2B81037C0C0B0003B42C3C4300743C3343F33C041E87008CCC280A32B89F0302C";
  defparam rom_dat0_2_0_11.INITVAL_12 = "0x200F00BCBF2F40C2B0A33B0CC3A03C03C8C3000F0880200023030002303030C080C0C83D03C220DC";
  defparam rom_dat0_2_0_11.INITVAL_13 = "0x0C8803C0C2040BC3003F3EC4C3080B3002000808088003CCC0000003F03C300083E0B1304B120030";
  defparam rom_dat0_2_0_11.INITVAL_14 = "0x018C636C960348008032000B704002258140840810C32010BC00028000CC0F070230700400630000";
  defparam rom_dat0_2_0_11.INITVAL_15 = "0x0000A000800D8C0010370DCC33280A100000C0F20ECA62ECC02000303043200B0320042A8540A040";
  defparam rom_dat0_2_0_11.INITVAL_16 = "0x03C413C8C2000323A0921003B10C06318C63C00226803000C000C210C8340C830098970CC800CC44";
  defparam rom_dat0_2_0_11.INITVAL_17 = "0x104102001000C003B84C0CCE82283A00C00008800203C1800302080300082000A1240020CDC0A801";
  defparam rom_dat0_2_0_11.INITVAL_18 = "0x0C0C0380003000C300033D0FF200003400E0000002CC0020C20004008808208000848003C0300CC0";
  defparam rom_dat0_2_0_11.INITVAL_19 = "0x3F008030042C48E2B8030380F06CFC300182E00C190E80F03300030200730000021408020FC38020";
  defparam rom_dat0_2_0_11.INITVAL_1A = "0x30CF03D0033AC03300FF1C03E0303C13C7F340300B84004C030C43020C233F0DF0DCB03FC330F0FF";
  defparam rom_dat0_2_0_11.INITVAL_1B = "0x36C331EC3336C331E8333B8333B833380EE0CCC3208EC2FC6C0B0030E80F380032F08C0F88F00C03";
  defparam rom_dat0_2_0_11.INITVAL_1C = "0x00CB3170E82883A08800380C31EC431E8D012C7C1C0B00F8000300F2000E0C03E000380D8331EC33";
  defparam rom_dat0_2_0_11.INITVAL_1D = "0x000F00FC00018E03C8023C0380000A0000220C303308F0C0CC33C012E41F0A41A02C28008A0000E0";
  defparam rom_dat0_2_0_11.INITVAL_1E = "0x000280043C008003202004000018CF308020C4C6318EC20C04300101C401030001000A294011A000";
  defparam rom_dat0_2_0_11.INITVAL_1F = "0x004002848E130C10282306C1E1086F28447004000F0103300E3D81C0C0333F0CC33C002107011009";
  defparam rom_dat0_2_0_11.INITVAL_20 = "0x20CF333C063C0030006E0F0883004000010200012D8EC1402C034000244002001008020001021055";
  defparam rom_dat0_2_0_11.INITVAL_21 = "0x14455104451500005000044551400300CC0000CC000000A0FC3BC043CC3C08C002D80308C3333801";
  defparam rom_dat0_2_0_11.INITVAL_22 = "0x15055054141145115045114551505404005054100540515405054540145000051044511044505455";
  defparam rom_dat0_2_0_11.INITVAL_23 = "0x15415154150541105415150551505415055150541105010040004100445514444150510440415444";
  defparam rom_dat0_2_0_11.INITVAL_24 = "0x05414154151541415414154141541411454154441545014445150541145115055154441544015410";
  defparam rom_dat0_2_0_11.INITVAL_25 = "0x00010000150400511040150441540005040000400144000040000151104415445054150541105415";
  defparam rom_dat0_2_0_11.INITVAL_26 = "0x00005154000000000001154050000510001050000144001010114050501111405040501400014000";
  defparam rom_dat0_2_0_11.INITVAL_27 = "0x00411000000000000000000000000014000140000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_11.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_11.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_11.INITVAL_2A = "0x000151FCEA2FCEA20015154400A8BF354400A8BF3FCEA20015100151FCEA2A8BF354400000000000";
  defparam rom_dat0_2_0_11.INITVAL_2B = "0x2A8BF35440054400A8BF3FCEA200151FCEA20015154400A8BF3A8BF35440000151FCEA2A8BF35440";
  defparam rom_dat0_2_0_11.INITVAL_2C = "0x0000000000000000005110044010401501414015000501045101404104150004111414100151FCEA";
  defparam rom_dat0_2_0_11.INITVAL_2D = "0x14CF0000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_11.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000008000000014000";
  defparam rom_dat0_2_0_11.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_11.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_11.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_11.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_11.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_11.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_11.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_11.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_11.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_11.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_11.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_11.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_11.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_11.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_11.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_11.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_11.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_11.OUTREG = "BYPASSED";
  defparam rom_dat0_2_0_11.RESETMODE = "SYNC";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:58226.9-58235.2" *)
  SP16K rom_dat0_2_0_12 (
    .AD({ builder_array_muxed0_12_RED_VOTER_wire, builder_array_muxed0_11_RED_VOTER_wire, builder_array_muxed0_10_RED_VOTER_wire, builder_array_muxed0_9_RED_VOTER_wire, builder_array_muxed0_8_RED_VOTER_wire, builder_array_muxed0_7_RED_VOTER_wire, builder_array_muxed0_6_RED_VOTER_wire, builder_array_muxed0_5_RED_VOTER_wire, builder_array_muxed0_4_RED_VOTER_wire, N_103_0_RED_VOTER_wire, builder_array_muxed0_2_RED_VOTER_wire, builder_array_muxed0_1_RED_VOTER_wire, builder_array_muxed0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire }),
    .CE(VCC_0_RED_VOTER_wire),
    .CLK(sys_clk),
    .CS({ VCC_0_RED_VOTER_wire, VCC_0_RED_VOTER_wire, VCC_0_RED_VOTER_wire }),
    .DI({ GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire }),
    .DO({ rom_dat0_2_0_12_DO, rom_dat0[25:24] }),
    .RST(GND_0_0_RED_VOTER_wire),
    .WE(GND_0_0_RED_VOTER_wire)
  );
  defparam rom_dat0_2_0_12.DATA_WIDTH = "X2";
  defparam rom_dat0_2_0_12.GSR = "ENABLED";
  defparam rom_dat0_2_0_12.INITVAL_00 = "0x0C005168AB0300101004074553E4581100000C020C80000830210000145A2BCF4154502A8AA00003";
  defparam rom_dat0_2_0_12.INITVAL_01 = "0x054110F40B0D01029C6437CFD14C341082004444340441C010084DE13C21360151E00E140071FCE7";
  defparam rom_dat0_2_0_12.INITVAL_02 = "0x33C140400226C5E154C121078124F30DCC43CCC43C01C370B435CD3184010185810C5C160C4048CC";
  defparam rom_dat0_2_0_12.INITVAL_03 = "0x110300440D14028000003241D0E04804050000C400CC80DCFE3AC00000C000000300000400800CFE";
  defparam rom_dat0_2_0_12.INITVAL_04 = "0x2003016855140E20602021C0401051188C001074144412A8FF08052060C00881100000020463C80D";
  defparam rom_dat0_2_0_12.INITVAL_05 = "0x08000000280082000088088500E0010002401403018220F8031308321409138310380405CC00546A";
  defparam rom_dat0_2_0_12.INITVAL_06 = "0x00028000003200115803040A002038008300540014804004002800320805140002C0302800510020";
  defparam rom_dat0_2_0_12.INITVAL_07 = "0x00003168A10801728004258031400F09C04080030009534803000023C01018025348030008300043";
  defparam rom_dat0_2_0_12.INITVAL_08 = "0x2800D340200800100030080F000800368A90803E100221F002044840201A24000100010001000C40";
  defparam rom_dat0_2_0_12.INITVAL_09 = "0x0001000022028031000C020251742000400008302080022400140001000C030000800D1A8AC20096";
  defparam rom_dat0_2_0_12.INITVAL_0A = "0x200390008914000300000001008CC0000080E000300352A81200079000891002C3E0003008215412";
  defparam rom_dat0_2_0_12.INITVAL_0B = "0x208632A000300833E03D01C9333C01210243C0D0034030000100010080C0000020F000300031A884";
  defparam rom_dat0_2_0_12.INITVAL_0C = "0x00020280000046A2FCC003000230CA0301401CFD07CC700C8D1C441310ED308D03E0310384F3F001";
  defparam rom_dat0_2_0_12.INITVAL_0D = "0x324A82B000024E9004C8000001000000860010CD070B00081E0841230000008C3000300008809003";
  defparam rom_dat0_2_0_12.INITVAL_0E = "0x220FD03080380390C8023780200C5014806108010880C0200011001300DA2AC20030440080C00001";
  defparam rom_dat0_2_0_12.INITVAL_0F = "0x040A9100501800208040040292C00205007008000381B104821040500C2210C00384020300801C27";
  defparam rom_dat0_2_0_12.INITVAL_10 = "0x2A84D30419100243C0020EC48088A73B8C3038840180023097148100780A124300147224C6008480";
  defparam rom_dat0_2_0_12.INITVAL_11 = "0x0280427C0C3501009C2025828200AA1100E080202D0A03200E38C463C002250C700029270160B080";
  defparam rom_dat0_2_0_12.INITVAL_12 = "0x000C80F4860380823020138812402C1244B24002200010000003801000300E0803808C0000801004";
  defparam rom_dat0_2_0_12.INITVAL_13 = "0x0C0070C0C03040C3803F0000E300103000320800000E002C80000C00000038000300392040E0B072";
  defparam rom_dat0_2_0_12.INITVAL_14 = "0x200151A8B6334000803000013080011589539C8200C000905E00002200433A0A8220300040008000";
  defparam rom_dat0_2_0_12.INITVAL_15 = "0x1C0000002007802000382B0823646202000000381C88F2284002002000801008C03000354553A853";
  defparam rom_dat0_2_0_12.INITVAL_16 = "0x0140D0C00001060000030800823C000546A2C000240372200300C000300002C34000C220C611C438";
  defparam rom_dat0_2_0_12.INITVAL_17 = "0x00C02040201500806CD1038B4104050008C044520846327056000C53005A0A41C030080583115408";
  defparam rom_dat0_2_0_12.INITVAL_18 = "0x1084C3200220002000080C00F00820300192081000C8030082080300C4031B4220A08C0040C154C2";
  defparam rom_dat0_2_0_12.INITVAL_19 = "0x240A10102001444000820002300000088100480811000230C2000B0010C20A00001452040100100C";
  defparam rom_dat0_2_0_12.INITVAL_1A = "0x00000300500000000000000C00000100C8000002090010005400C41004013041411C001C40100000";
  defparam rom_dat0_2_0_12.INITVAL_1B = "0x00C0300C0300C0300C030C0030C003000C000C03020B030C0C0005000000300080602C0000C00000";
  defparam rom_dat0_2_0_12.INITVAL_1C = "0x308001400825C000C80003C422045220093008B81C030000002C01000008300400002C0400300C03";
  defparam rom_dat0_2_0_12.INITVAL_1D = "0x2100110008100000001400030000C000004038000000000000000091441302412028280002801000";
  defparam rom_dat0_2_0_12.INITVAL_1E = "0x010031B02C0040000820000470100300C06068BF3002C10C2C300103C83303008000073FCD330C00";
  defparam rom_dat0_2_0_12.INITVAL_1F = "0x1480002090010032180B00055344E00809400402100133342E0180900024000D000C013309231041";
  defparam rom_dat0_2_0_12.INITVAL_20 = "0x00030000000401001401030401004000403008400146C3800001C002040001000000000081331015";
  defparam rom_dat0_2_0_12.INITVAL_21 = "0x10810210CA1005514415080732C080008040000100000080000042000C2000C10014000503012481";
  defparam rom_dat0_2_0_12.INITVAL_22 = "0x1307303031304F30F00C01C301F09C180093908026C66034001006C204B0000120C842104C90B096";
  defparam rom_dat0_2_0_12.INITVAL_23 = "0x2C4821680F03C1000C313F0CE1F0783707C3F08401430100200082000CD41008014C62074402C007";
  defparam rom_dat0_2_0_12.INITVAL_24 = "0x1900C1C00C0C00C1C41C1100C1101C1F00C05CC627C39244970900C01C3F03082110C7110C02C480";
  defparam rom_dat0_2_0_12.INITVAL_25 = "0x02CC2348870846C100A6310B4150930FCC431CC1070C3044F300417000CC21C0D0FC2F07C343C026";
  defparam rom_dat0_2_0_12.INITVAL_26 = "0x0000000000000000CC320101021453344502481514C551245422C400B4201EC4409CB4284550F454";
  defparam rom_dat0_2_0_12.INITVAL_27 = "0x00C0100000000000000000000008AA28455140000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_12.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_12.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_12.INITVAL_2A = "0x06C243C48E1C48E16C24390DB03871290DB038712C48E16C2436C243C48E13871290DB0000000000";
  defparam rom_dat0_2_0_12.INITVAL_2B = "0x13871290DB090DB038712C48E16C243C48E16C24390DB0387123871290DB06C243C48E13871290DB";
  defparam rom_dat0_2_0_12.INITVAL_2C = "0x00000000000000000000004940640139040120120805000032228251585C040432183826C243C48E";
  defparam rom_dat0_2_0_12.INITVAL_2D = "0x0CCF0000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_12.INITVAL_2E = "0x0000000000000000000000000000000000000000000000000000000000000000000800000000C000";
  defparam rom_dat0_2_0_12.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_12.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_12.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_12.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_12.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_12.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_12.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_12.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_12.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_12.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_12.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_12.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_12.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_12.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_12.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_12.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_12.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_12.OUTREG = "BYPASSED";
  defparam rom_dat0_2_0_12.RESETMODE = "SYNC";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:58145.9-58154.2" *)
  SP16K rom_dat0_2_0_13 (
    .AD({ builder_array_muxed0_12_RED_VOTER_wire, builder_array_muxed0_11_RED_VOTER_wire, builder_array_muxed0_10_RED_VOTER_wire, builder_array_muxed0_9_RED_VOTER_wire, builder_array_muxed0_8_RED_VOTER_wire, builder_array_muxed0_7_RED_VOTER_wire, builder_array_muxed0_6_RED_VOTER_wire, builder_array_muxed0_5_RED_VOTER_wire, builder_array_muxed0_4_RED_VOTER_wire, N_103_0_RED_VOTER_wire, builder_array_muxed0_2_RED_VOTER_wire, builder_array_muxed0_1_RED_VOTER_wire, builder_array_muxed0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire }),
    .CE(VCC_0_RED_VOTER_wire),
    .CLK(sys_clk),
    .CS({ VCC_0_RED_VOTER_wire, VCC_0_RED_VOTER_wire, VCC_0_RED_VOTER_wire }),
    .DI({ GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire }),
    .DO({ rom_dat0_2_0_13_DO, rom_dat0[27:26] }),
    .RST(GND_0_0_RED_VOTER_wire),
    .WE(GND_0_0_RED_VOTER_wire)
  );
  defparam rom_dat0_2_0_13.DATA_WIDTH = "X2";
  defparam rom_dat0_2_0_13.GSR = "ENABLED";
  defparam rom_dat0_2_0_13.INITVAL_00 = "0x0000000003030100001404000000000700308C0304C000080011010000000000F3FCFF3FCFF00002";
  defparam rom_dat0_2_0_13.INITVAL_01 = "0x000000F0010C000014402FC3F000300040100000100000C000040ED03C23120D414008100000F047";
  defparam rom_dat0_2_0_13.INITVAL_02 = "0x33800000032F84C330000007D03CF30CCC03C0C00C44C130B030CB33004004C0900404000000000C";
  defparam rom_dat0_2_0_13.INITVAL_03 = "0x040A9330000004800800110022E01000010000000400704000008C20008000033380000400C00CBE";
  defparam rom_dat0_2_0_13.INITVAL_04 = "0x0403000000040200C0C031800000000141000030000040000009C9004CC00D000000002300E18CCC";
  defparam rom_dat0_2_0_13.INITVAL_05 = "0x0000F0000C000300100C00C300E000200080140331CDA05000030A73043D03C10034000004000000";
  defparam rom_dat0_2_0_13.INITVAL_06 = "0x0003C00000300000080D0C0C00000800C100000000C0C000003C0032000000000000003800000033";
  defparam rom_dat0_2_0_13.INITVAL_07 = "0x010000000A00020000000FC00080070880838000000001800100003240303400034003000C010004";
  defparam rom_dat0_2_0_13.INITVAL_08 = "0x000031803004008000200009000C00000010000000000340000C0C30300004000300080000008840";
  defparam rom_dat0_2_0_13.INITVAL_09 = "0x004000003A02C022000800000038000000000C5004C0100C002C0020100802C000C0000000800000";
  defparam rom_dat0_2_0_13.INITVAL_0A = "0x0004000003200000400400030004C0000040800000000000A000800000033C024380003000000060";
  defparam rom_dat0_2_0_13.INITVAL_0B = "0x2848114009040821B0D7334E3134100000C08470318A910005000200005000C00080003008000018";
  defparam rom_dat0_2_0_13.INITVAL_0C = "0x01000080000040000015134C02104E0340A0000118008118A52440300C4204C501C010010C4114E1";
  defparam rom_dat0_2_0_13.INITVAL_0D = "0x0200003C0000003300D800030000C0094C8024631400000019060803401000C4514034000010F412";
  defparam rom_dat0_2_0_13.INITVAL_0E = "0x330FD03010140330408133800000551580620C490442C22008200033000000C20030800000C00082";
  defparam rom_dat0_2_0_13.INITVAL_0F = "0x000A6100F0000C000010000033C40402001008400308B2C00220C300946930400000470000C08C93";
  defparam rom_dat0_2_0_13.INITVAL_10 = "0x24C0C20832200C33C0C00C00800800334C103098004000380F0C8CC0380C014051547030C102C020";
  defparam rom_dat0_2_0_13.INITVAL_11 = "0x244000AC04330003000004C00000810101504838360961180D3140B3C0002E0C3000003701301000";
  defparam rom_dat0_2_0_13.INITVAL_12 = "0x000E00B88A324040F000034470000C03C4000008300030000003000000300CC8E34844228200A004";
  defparam rom_dat0_2_0_13.INITVAL_13 = "0x0C0033F0C03000C3003B0000F300003000310C00000F003CC0000F000000300003A0321000000030";
  defparam rom_dat0_2_0_13.INITVAL_14 = "0x00000000A303000080330000300000000000388300C000000C00003204200000800CFC0000000000";
  defparam rom_dat0_2_0_13.INITVAL_15 = "0x0000120815110200C048020043DC3303C000007D04005154003100000020000CC030C00545515460";
  defparam rom_dat0_2_0_13.INITVAL_16 = "0x02008000300043000003048B411015154551F000100330008000C400DC0001812000C010C8008032";
  defparam rom_dat0_2_0_13.INITVAL_17 = "0x004010C4020000C044800146008020040C0200010003430803000003900E0A04C0308A00C5C0C00C";
  defparam rom_dat0_2_0_13.INITVAL_18 = "0x00C4C33003300030000C0C00F000303002C3000400C100300000818044030B0200E0880080830CC3";
  defparam rom_dat0_2_0_13.INITVAL_19 = "0x20001010000000000010000132C00000400000002300003C00000B0000000000000003000300100C";
  defparam rom_dat0_2_0_13.INITVAL_1A = "0x00000300000000000000000C00000000C0000000000410400001C00000803000000C000C00000000";
  defparam rom_dat0_2_0_13.INITVAL_1B = "0x00C0300C0300C0300C030C0030C003000F000C00000303400C0C00000000000000303C0000C00000";
  defparam rom_dat0_2_0_13.INITVAL_1C = "0x3000014008284010840003840100D0100001007010030000000C00000001300000000C0800300C03";
  defparam rom_dat0_2_0_13.INITVAL_1D = "0x31000000000003000000000B0000C80000003C20000800800020000014120141602C180002C00012";
  defparam rom_dat0_2_0_13.INITVAL_1E = "0x000030F02800040000000400200001000040000005454208083002024C22030000C0000001405808";
  defparam rom_dat0_2_0_13.INITVAL_1F = "0x00000034C00100002C3100000308C003400008020001111004000D800030000C200C00320310000C";
  defparam rom_dat0_2_0_13.INITVAL_20 = "0x00C92088002C0200300A010B03008100030200000001414024020001008002003000000082033040";
  defparam rom_dat0_2_0_13.INITVAL_21 = "0x20C740500C310FF31C3F080F7300C03CC880CC00088220C0E328C000BCF900420028030881033802";
  defparam rom_dat0_2_0_13.INITVAL_22 = "0x000400C001024301307101C44030C01C04800C1024047304271640C21030020921C4A0344090FC17";
  defparam rom_dat0_2_0_13.INITVAL_23 = "0x3E4972741304C1104C053301F130FF0B08C3308431070008200000020067228C03ACB30441010004";
  defparam rom_dat0_2_0_13.INITVAL_24 = "0x3041C0141C0141C0182C1341C1341C1300C3C0C534C33348C70805C1D018170D0260C4060C83E498";
  defparam rom_dat0_2_0_13.INITVAL_25 = "0x2A052100870B4C42148C120A8014323FCCC23CC30F0C30CCF300C27110CC1DC4E00C0300C0C21434";
  defparam rom_dat0_2_0_13.INITVAL_26 = "0x000000000000000000030303B03CF20CCF11803F3CC3F304FC268C51AC24328C6090AC10CFF0ECFC";
  defparam rom_dat0_2_0_13.INITVAL_27 = "0x00C32000000000000000000000000000000000500000200000000000000000000000000000000000";
  defparam rom_dat0_2_0_13.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_13.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_13.INITVAL_2A = "0x0E06D01C923B438148C7248C72B438148C72B4381B438148C72E06D01C9231C923E06D0000000000";
  defparam rom_dat0_2_0_13.INITVAL_2B = "0x31C923E06D048C72B4381B438148C72B438148C7248C72B43811C923E06D0E06D01C9231C923E06D";
  defparam rom_dat0_2_0_13.INITVAL_2C = "0x00000000000000000010134103444D01044100100C09012042020272505D0C8C133C2C0E06D01C92";
  defparam rom_dat0_2_0_13.INITVAL_2D = "0x00CF0000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_13.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000004000000000000";
  defparam rom_dat0_2_0_13.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_13.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_13.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_13.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_13.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_13.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_13.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_13.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_13.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_13.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_13.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_13.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_13.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_13.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_13.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_13.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_13.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_13.OUTREG = "BYPASSED";
  defparam rom_dat0_2_0_13.RESETMODE = "SYNC";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:58064.9-58073.2" *)
  SP16K rom_dat0_2_0_14 (
    .AD({ builder_array_muxed0_12_RED_VOTER_wire, builder_array_muxed0_11_RED_VOTER_wire, builder_array_muxed0_10_RED_VOTER_wire, builder_array_muxed0_9_RED_VOTER_wire, builder_array_muxed0_8_RED_VOTER_wire, builder_array_muxed0_7_RED_VOTER_wire, builder_array_muxed0_6_RED_VOTER_wire, builder_array_muxed0_5_RED_VOTER_wire, builder_array_muxed0_4_RED_VOTER_wire, N_103_0_RED_VOTER_wire, builder_array_muxed0_2_RED_VOTER_wire, builder_array_muxed0_1_RED_VOTER_wire, builder_array_muxed0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire }),
    .CE(VCC_0_RED_VOTER_wire),
    .CLK(sys_clk),
    .CS({ VCC_0_RED_VOTER_wire, VCC_0_RED_VOTER_wire, VCC_0_RED_VOTER_wire }),
    .DI({ GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire }),
    .DO({ rom_dat0_2_0_14_DO, rom_dat0[29:28] }),
    .RST(GND_0_0_RED_VOTER_wire),
    .WE(GND_0_0_RED_VOTER_wire)
  );
  defparam rom_dat0_2_0_14.DATA_WIDTH = "X2";
  defparam rom_dat0_2_0_14.GSR = "ENABLED";
  defparam rom_dat0_2_0_14.INITVAL_00 = "0x0000000003030000000000000000000300130C0315C0004477334C0000000000B3FCFF3FCFF00000";
  defparam rom_dat0_2_0_14.INITVAL_01 = "0x00000070002C000000002FCFE0003000C000C000000000C0010CCFC03C33030C0030083000003042";
  defparam rom_dat0_2_0_14.INITVAL_02 = "0x33C000002333C8C33000000CC03CFB0CCD03C4C01C44C330F0100F03000000C0F00000000200088C";
  defparam rom_dat0_2_0_14.INITVAL_03 = "0x0C0F83300800008008C00002A0B0D00000C00080300070545515C8200040000F01C8000C00C00CFD";
  defparam rom_dat0_2_0_14.INITVAL_04 = "0x0001000000000100F0830000000000048400003000005154550400304CCD0408000000320470C4C4";
  defparam rom_dat0_2_0_14.INITVAL_05 = "0x0000F0000C000300000C00000000040000C00003318D304C0003040300180340001000020C000000";
  defparam rom_dat0_2_0_14.INITVAL_06 = "0x0403C000432000000C0B0C09000004044300000100C0C00000140033000000000040001400000033";
  defparam rom_dat0_2_0_14.INITVAL_07 = "0x020000000100020000000C8010804B0D40C34003000001400300003140331400014003000C210059";
  defparam rom_dat0_2_0_14.INITVAL_08 = "0x000032C0300C00F00000000F0000000000F00010000003F00F0C0C3030000C0001000F0002000C40";
  defparam rom_dat0_2_0_14.INITVAL_09 = "0x0080000030034030000800000004000C00000C4030C0300C001C0033000C03C000C0000002C00000";
  defparam rom_dat0_2_0_14.INITVAL_0A = "0x0000000003280033000D0000000C00010000F00010000000D000400000033003C3F0001000000010";
  defparam rom_dat0_2_0_14.INITVAL_0B = "0x0000000000000003303C30C3030C7131C18184F3300033000E00030000E000C000E0003000000024";
  defparam rom_dat0_2_0_14.INITVAL_0C = "0x0000000000000000000003040000050301A000000801804CF534C0200CC000C500D0310200033000";
  defparam rom_dat0_2_0_14.INITVAL_0D = "0x010000300000003300C800020000800A8D4034F3050000000A0208030030004C200430000440F030";
  defparam rom_dat0_2_0_14.INITVAL_0E = "0x1103C00010000020404000400000000040310C091986D2700C100032000000C10030400040C00003";
  defparam rom_dat0_2_0_14.INITVAL_0F = "0x00071100F00004000010000013C00005000004800308C20002008203003330C003008B0000400C00";
  defparam rom_dat0_2_0_14.INITVAL_10 = "0x1CC0C10C22100C31C0E00C00400400338C203074000000300F0840002400000000003130C303C030";
  defparam rom_dat0_2_0_14.INITVAL_11 = "0x200010FC0C330201082000C00000400105A08879380622684E3081B0C040150C2000303703301000";
  defparam rom_dat0_2_0_14.INITVAL_12 = "0x000E10FCCF33C0C0F000030030000C0000001000300020000003000000300C80E398892286009005";
  defparam rom_dat0_2_0_14.INITVAL_13 = "0x0C003330003000C3003F0000F000000000300C00000F003CC0000F000000300003840224C330C030";
  defparam rom_dat0_2_0_14.INITVAL_14 = "0x00000000F3000000000000001000080000003CC300C000000C00003100100000400CFC0000000000";
  defparam rom_dat0_2_0_14.INITVAL_15 = "0x0D81308031030300000C030000CC3300C000000C00000000003200000020000CC030800000000030";
  defparam rom_dat0_2_0_14.INITVAL_16 = "0x070000C00000030000030200000000000000F00020033000C200C0000C0000800000C0000C00CCFE";
  defparam rom_dat0_2_0_14.INITVAL_17 = "0x01802084022000C00080000100401004040100010003430403000003400D0500C0306400C4C0C02C";
  defparam rom_dat0_2_0_14.INITVAL_18 = "0x00C0C33003300030000C0C00F000303001C3000800C200300000808000030B0000E0880080430C0B";
  defparam rom_dat0_2_0_14.INITVAL_19 = "0x01001010000000000020000031000000C00008083200003C0000000010000000000003000300000C";
  defparam rom_dat0_2_0_14.INITVAL_1A = "0x000000000000000000000000000C0000C800C000080000C0000080C000C03000000C000C00000000";
  defparam rom_dat0_2_0_14.INITVAL_1B = "0x00C0000C0000C0000C000C0000C000000F000000000303000C0C00000000000000303C0000C00000";
  defparam rom_dat0_2_0_14.INITVAL_1C = "0x300001400B280030800003C00000C0000030003030030000000C0000003030000000C00800000C00";
  defparam rom_dat0_2_0_14.INITVAL_1D = "0x3300000000000300000000030000000000003030000C00C000300000041100412024080002C00020";
  defparam rom_dat0_2_0_14.INITVAL_1E = "0x000030E030000C0000000C0C00000300C00000000003C00000300303C00003000000000000000C0C";
  defparam rom_dat0_2_0_14.INITVAL_1F = "0x0040003CC0030001200300000044800004403000000D13142C00004100F0000C000C0E0208120000";
  defparam rom_dat0_2_0_14.INITVAL_20 = "0x07C82008002F4640F00A000B037490000F310000000343403403400000C002001000080201000000";
  defparam rom_dat0_2_0_14.INITVAL_21 = "0x388EE2C8CB2B0FF2B8BF038AA280403CC990CC00398661C0E320C430BCF813024028530880037812";
  defparam rom_dat0_2_0_14.INITVAL_22 = "0x270AF0B832328A32A0EE228BC2A0EC288CE2A8300B8AE2B83E2F8900E840030E328C43208820A8EE";
  defparam rom_dat0_2_0_14.INITVAL_23 = "0x2B8EE3A82A0A83A2A43A2A0EA2A06F3D0A82A0EE2A8D33FC8F3E4FF38CBA2288C2E8A20B8BB2EC0A";
  defparam rom_dat0_2_0_14.INITVAL_24 = "0x2AC342E8243EC342EC342AC342AC242A8C42A88B2A82D2A8E90E8B43A827290BB2A84A2A84F2B8EF";
  defparam rom_dat0_2_0_14.INITVAL_25 = "0x3FCB03FC2C00CBB230BB2E01A2B821354681A4AA0A86A288592A83A330880A8CA0E83A0E8361EC2B";
  defparam rom_dat0_2_0_14.INITVAL_26 = "0x0000000000000000CC322A02E33CF93ACF22A83F3F8FF308880B48F2D80A2F4800ECD834CFF39CFC";
  defparam rom_dat0_2_0_14.INITVAL_27 = "0x0082000000000000000000000010000100001405168AA28000000000000000000000000000000000";
  defparam rom_dat0_2_0_14.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_14.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_14.INITVAL_2A = "0x16C1B06C1B0C4B12C4B1290E4390E43C4B12C4B1290E4390E43384E1384E16C1B06C1B0000000000";
  defparam rom_dat0_2_0_14.INITVAL_2B = "0x3C4B12C4B126C1B06C1B0384E1384E16C1B06C1B0384E1384E190E4390E43C4B12C4B12384E1384E";
  defparam rom_dat0_2_0_14.INITVAL_2C = "0x000001545515455140B2328E82B88A3F0AC2902B088B2228B313C0A2ACA700CB020808090E4390E4";
  defparam rom_dat0_2_0_14.INITVAL_2D = "0x04CF0000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_14.INITVAL_2E = "0x0000000000000000000000000000000000000000000000000000000000000000000C400000004000";
  defparam rom_dat0_2_0_14.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_14.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_14.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_14.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_14.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_14.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_14.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_14.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_14.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_14.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_14.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_14.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_14.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_14.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_14.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_14.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_14.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_14.OUTREG = "BYPASSED";
  defparam rom_dat0_2_0_14.RESETMODE = "SYNC";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57983.9-57992.2" *)
  SP16K rom_dat0_2_0_15 (
    .AD({ builder_array_muxed0_12_RED_VOTER_wire, builder_array_muxed0_11_RED_VOTER_wire, builder_array_muxed0_10_RED_VOTER_wire, builder_array_muxed0_9_RED_VOTER_wire, builder_array_muxed0_8_RED_VOTER_wire, builder_array_muxed0_7_RED_VOTER_wire, builder_array_muxed0_6_RED_VOTER_wire, builder_array_muxed0_5_RED_VOTER_wire, builder_array_muxed0_4_RED_VOTER_wire, N_103_0_RED_VOTER_wire, builder_array_muxed0_2_RED_VOTER_wire, builder_array_muxed0_1_RED_VOTER_wire, builder_array_muxed0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire }),
    .CE(VCC_0_RED_VOTER_wire),
    .CLK(sys_clk),
    .CS({ VCC_0_RED_VOTER_wire, VCC_0_RED_VOTER_wire, VCC_0_RED_VOTER_wire }),
    .DI({ GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire }),
    .DO({ rom_dat0_2_0_15_DO, rom_dat0[31:30] }),
    .RST(GND_0_0_RED_VOTER_wire),
    .WE(GND_0_0_RED_VOTER_wire)
  );
  defparam rom_dat0_2_0_15.DATA_WIDTH = "X2";
  defparam rom_dat0_2_0_15.GSR = "ENABLED";
  defparam rom_dat0_2_0_15.INITVAL_00 = "0x0000000007030000001000000000000300108C0100C00080303300000000000033FCFF3FCFF00000";
  defparam rom_dat0_2_0_15.INITVAL_01 = "0x000000F0003C000000003FCFF0003000C000C000000000C0000CCFC03C33030C0000003000003000";
  defparam rom_dat0_2_0_15.INITVAL_02 = "0x33C000003333CCC33000000CC03CFF0CCF03CCC03CCCC330F0300F03000000C0F000000003000CCC";
  defparam rom_dat0_2_0_15.INITVAL_03 = "0x0E0F03B8022A800004C000000030040800C288A23044000000000C20000000021000000000C00CBF";
  defparam rom_dat0_2_0_15.INITVAL_04 = "0x0001000000040200F05300C000000000C00000300000000000000030040C0004000000330030C0C0";
  defparam rom_dat0_2_0_15.INITVAL_05 = "0x0000F0000C000300000C00410050041000007C03314D705C10030503001403410014000100000000";
  defparam rom_dat0_2_0_15.INITVAL_06 = "0x0403C030233000000C000C01000008048000000100C0C00000280033000000000040002800000033";
  defparam rom_dat0_2_0_15.INITVAL_07 = "0x010000000100010000000C400040070C40434001000000400100003040330400004001000C010001";
  defparam rom_dat0_2_0_15.INITVAL_08 = "0x00003140300C00D00010000D0004000000500010000003500D0C0C3030000C0001000D0001000C40";
  defparam rom_dat0_2_0_15.INITVAL_09 = "0x000000003603C032000000000014000000000C6038C0320C00140031000003400000000001400040";
  defparam rom_dat0_2_0_15.INITVAL_0A = "0x0000000003080033000E0000000C80000000D00000000000100000000003080303D0000000000050";
  defparam rom_dat0_2_0_15.INITVAL_0B = "0x300C03C003300300200820020200202080808000200033000E00010000E0004000E0001000000004";
  defparam rom_dat0_2_0_15.INITVAL_0C = "0x00000040000000000000030001000A03010000000000000CDF1C80200401004F017003030CC000C0";
  defparam rom_dat0_2_0_15.INITVAL_0D = "0x020000300000003300CC00030000C0030DC03433050000000C00000300100040000030000000F031";
  defparam rom_dat0_2_0_15.INITVAL_0E = "0x1103C00000000030000000000000000080320C010000C03000300030000000C20000C00040C04000";
  defparam rom_dat0_2_0_15.INITVAL_0F = "0x000B3300E0000C000020000003C0000300000800130CC3C00300C340000330C00000CF0000C00C00";
  defparam rom_dat0_2_0_15.INITVAL_10 = "0x28C0C10831310831C0D008008008C0334C10309C0000007C0F048CC0180C000000003330C103D010";
  defparam rom_dat0_2_0_15.INITVAL_11 = "0x000000CC0C300342041000C04000800100000030390800000C3000F1C040270C1000603703301000";
  defparam rom_dat0_2_0_15.INITVAL_12 = "0x100C00FCCF33C0C0F000030030000C0000000000300030000003000000300CC4C200000000001004";
  defparam rom_dat0_2_0_15.INITVAL_13 = "0x0C003330003000C3003F0000F000000000300C04000F003CC0000F010000300003000300C330C030";
  defparam rom_dat0_2_0_15.INITVAL_14 = "0x00000000F3000000400100013000000000003CC300C000000C00003200000000800CFC0000000000";
  defparam rom_dat0_2_0_15.INITVAL_15 = "0x0C00300030030700000C030000CC3300C000000C00000000003000000000000CC030000000000030";
  defparam rom_dat0_2_0_15.INITVAL_16 = "0x034010800000035140030000000000000000F00004037000C200C0000C0000C00000C0000C00CCFC";
  defparam rom_dat0_2_0_15.INITVAL_17 = "0x00C0308C030008C000C00000011004000C0000400003030003000003000C0000C0300000C0D0D00C";
  defparam rom_dat0_2_0_15.INITVAL_18 = "0x00C0C37003300070000C0C00F000303002D2003C00CF00300400C7C000031F0300F4CC00C0C30C03";
  defparam rom_dat0_2_0_15.INITVAL_19 = "0x00004000000000000400000030000010C00010003000003C0000000000000000000003000300000C";
  defparam rom_dat0_2_0_15.INITVAL_1A = "0x000000000001400100010000400C0400CC01C0000C4000C00004C0C000D03404400C000C00000001";
  defparam rom_dat0_2_0_15.INITVAL_1B = "0x00C0000C0000C0000C000C0000C000000F000001000303140C0C0000000100000020380004D00000";
  defparam rom_dat0_2_0_15.INITVAL_1C = "0x300001400B2C8030C80003C80040E0040072000038000004080E02A208B0380AA028C40C00000C00";
  defparam rom_dat0_2_0_15.INITVAL_1D = "0x3300000400000300000004030000C00000003030000C00C00030000004130041202C080002C00032";
  defparam rom_dat0_2_0_15.INITVAL_1E = "0x000030F028000C000000080CE0000200C000000000020308003002020C2003000000000000000C0C";
  defparam rom_dat0_2_0_15.INITVAL_1F = "0x0080003CC0030002382000000288C4120AA030002A0E20282C1108A280F0000E822CAE220A020008";
  defparam rom_dat0_2_0_15.INITVAL_20 = "0x00C0000000070000F0000003013000000F3200000003838038038000008002002000000002222080";
  defparam rom_dat0_2_0_15.INITVAL_21 = "0x1005415041110001140000055140C02CC0008800300000C0C20040302CB000000040030000013000";
  defparam rom_dat0_2_0_15.INITVAL_22 = "0x15055050100145115055004541501404001150500545511404054540145001040140511444105055";
  defparam rom_dat0_2_0_15.INITVAL_23 = "0x15015154150541104415150551505015054150441145000400004001045511444154510545110405";
  defparam rom_dat0_2_0_15.INITVAL_24 = "0x15414154141541415414114141141415044154451541514415050541541515011150451504015010";
  defparam rom_dat0_2_0_15.INITVAL_25 = "0x00450000450100501440140041545115444104010404004451004151104415445014050140415415";
  defparam rom_dat0_2_0_15.INITVAL_26 = "0x00000000000000004411010150000014001144000040001054040451040404045044041400005000";
  defparam rom_dat0_2_0_15.INITVAL_27 = "0x00411000000000000000000000000014000140000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_15.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_15.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_15.INITVAL_2A = "0x1E0781E0781E0781E0781E0781E0781B42D0B42D0B42D0B42D0B42D0B42D0B42D0B42D0000000000";
  defparam rom_dat0_2_0_15.INITVAL_2B = "0x21C8721C8721C8721C8721C8721C87248D2348D2348D2348D2348D2348D2348D2348D23E0781E078";
  defparam rom_dat0_2_0_15.INITVAL_2C = "0x000000000000000000101105411444150041101100050100501040514455004010101011C8721C87";
  defparam rom_dat0_2_0_15.INITVAL_2D = "0x04CF0000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_15.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000004000";
  defparam rom_dat0_2_0_15.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_15.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_15.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_15.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_15.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_15.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_15.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_15.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_15.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_15.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_15.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_15.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_15.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_15.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_15.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_15.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_15.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_15.OUTREG = "BYPASSED";
  defparam rom_dat0_2_0_15.RESETMODE = "SYNC";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:59036.9-59045.2" *)
  SP16K rom_dat0_2_0_2 (
    .AD({ builder_array_muxed0_12_RED_VOTER_wire, builder_array_muxed0_11_RED_VOTER_wire, builder_array_muxed0_10_RED_VOTER_wire, builder_array_muxed0_9_RED_VOTER_wire, builder_array_muxed0_8_RED_VOTER_wire, builder_array_muxed0_7_RED_VOTER_wire, builder_array_muxed0_6_RED_VOTER_wire, builder_array_muxed0_5_RED_VOTER_wire, builder_array_muxed0_4_RED_VOTER_wire, N_103_0_RED_VOTER_wire, builder_array_muxed0_2_RED_VOTER_wire, builder_array_muxed0_1_RED_VOTER_wire, builder_array_muxed0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire }),
    .CE(VCC_0_RED_VOTER_wire),
    .CLK(sys_clk),
    .CS({ VCC_0_RED_VOTER_wire, VCC_0_RED_VOTER_wire, VCC_0_RED_VOTER_wire }),
    .DI({ GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire }),
    .DO({ rom_dat0_2_0_2_DO, rom_dat0[5:4] }),
    .RST(GND_0_0_RED_VOTER_wire),
    .WE(GND_0_0_RED_VOTER_wire)
  );
  defparam rom_dat0_2_0_2.DATA_WIDTH = "X2";
  defparam rom_dat0_2_0_2.GSR = "ENABLED";
  defparam rom_dat0_2_0_2.INITVAL_00 = "0x2400000009350A321455158AA2A8AB3D06A378691585825457154D000000000092A8AA2A8AA15456";
  defparam rom_dat0_2_0_2.INITVAL_01 = "0x2A8761988A268381D459294962881D298220A899190DA2706609866354261A4A626459290BE1589A";
  defparam rom_dat0_2_0_2.INITVAL_02 = "0x088AA1E462268A62A4A3224963D8582242D1484D248A4290992A45918C861B8F6248A83A4A90D894";
  defparam rom_dat0_2_0_2.INITVAL_03 = "0x2A4692286A2A8A9154D7260EA2A4A72145D2986E384793A8AA2A47A14085150F6278A916C662A496";
  defparam rom_dat0_2_0_2.INITVAL_04 = "0x0BCED2A8AA274863649E258D314C540989B14C531402400000198A22A8791989535C5026C4A2A8AA";
  defparam rom_dat0_2_0_2.INITVAL_05 = "0x1649A0B468168661A0692585C094D91C06A1D06D264A6198FE164991346616853364761647000000";
  defparam rom_dat0_2_0_2.INITVAL_06 = "0x378291149719000008592949602025374E62A8BD2B48A1240216CE92640000814284261546A2F89A";
  defparam rom_dat0_2_0_2.INITVAL_07 = "0x12449000093842A29419264E6170A53A4D9278121484027812294192786B2749027812294461E849";
  defparam rom_dat0_2_0_2.INITVAL_08 = "0x29419278690BC59384250949E04852100093842A2506619C993989A1646A29455250993842509878";
  defparam rom_dat0_2_0_2.INITVAL_09 = "0x048A5064993A8561E04912490024E10A8512649E278D61E855254821E049124E10942400027210AA";
  defparam rom_dat0_2_0_2.INITVAL_0A = "0x210AA14499278A72945938C25098783244919C84250900009E048AA144992786919C84250990009E";
  defparam rom_dat0_2_0_2.INITVAL_0B = "0x1785E154F917C9E19C9A1E49E1E49E1E4E72786F368A925459384250949E0485219C842509900027";
  defparam rom_dat0_2_0_2.INITVAL_0C = "0x31421294281240000000064861E4953E495168AA268B62E4A526846158621785F29C993A87A1985E";
  defparam rom_dat0_2_0_2.INITVAL_0D = "0x1400309825128A926C9A0E063374851A8A51E86E194B607C5A188B6258660587829C65214991A466";
  defparam rom_dat0_2_0_2.INITVAL_0E = "0x2645A19C61190D93889215826258AA2A0B90E8653B8E72E84B12C72248400248E12C4B1C8F52D0A6";
  defparam rom_dat0_2_0_2.INITVAL_0F = "0x0A42917CA51548C1AC2832C522584909C72250BD3908929456134E5264A625836244563D835394A5";
  defparam rom_dat0_2_0_2.INITVAL_10 = "0x08824248621FC82250A50A8221208212852254271C8F52D8090908A12038090400001A224242B025";
  defparam rom_dat0_2_0_2.INITVAL_11 = "0x0982F0A44A1242F2886528849124220D4E2290E32A4280E0E61A07A250A509C723D4E02942212449";
  defparam rom_dat0_2_0_2.INITVAL_12 = "0x3A8672986619849184F62989935475124492644924C45358B209859320991687A2B093280E9124D7";
  defparam rom_dat0_2_0_2.INITVAL_13 = "0x148A92685A12406190992D84616090198A12486E09CA62E494264A63A03D1A49A19C9A0E8661989A";
  defparam rom_dat0_2_0_2.INITVAL_14 = "0x04000000AA15C951945615455254562A8AA298A60448A24406150A90E42A2A8612E49A1241009056";
  defparam rom_dat0_2_0_2.INITVAL_15 = "0x2949A164A61A4E52906B1ECE616866168460D09615455154552685612462154672DC902A8AA2A899";
  defparam rom_dat0_2_0_2.INITVAL_16 = "0x0644B094A7294573F841198661904000000068532EC6D2949616449098650986E1544619455168A9";
  defparam rom_dat0_2_0_2.INITVAL_17 = "0x118521989615C7B2649D3986D3BC6F194A525CE6194590D85527C95194563A455014991549919499";
  defparam rom_dat0_2_0_2.INITVAL_18 = "0x128A61E41A2506E2502B360F5258A51886B2946A134A9164652586A164563AC691A4992585A25866";
  defparam rom_dat0_2_0_2.INITVAL_19 = "0x2645E16491000133FC661ACAD2BCFD3586A278592E4AE2D8EB2B8A62A4EB2A4552A8A924425264A6";
  defparam rom_dat0_2_0_2.INITVAL_1A = "0x354F51D45B3FC573547F1D47D174FD17CBF3946519C9619CFF1D8AB354B51FCF73F4F5174751F4FF";
  defparam rom_dat0_2_0_2.INITVAL_1B = "0x3D0353D0353D0353D03533435334353486D0D4D13ECDD1B4753B4531D42B1DC64028592FCD715C57";
  defparam rom_dat0_2_0_2.INITVAL_1C = "0x1D8221E087394C21A4D5398771D49F1D49E1DC5B274992FC5D2A88A258BD2A82A168F72B4353D035";
  defparam rom_dat0_2_0_2.INITVAL_1D = "0x264B51FC5A100252CC573D49517C891546A2D8E52349B1948D26C64024720A47917825168B619429";
  defparam rom_dat0_2_0_2.INITVAL_1E = "0x37469264651ACA508865094991B8D2258641000000027254EB1546C2785E1D4780945A2A8AA2A499";
  defparam rom_dat0_2_0_2.INITVAL_1F = "0x2A4D529890020D7264E530000278BF3DC86378560A4E21E4EB3FC781B4E62A44A264AE1E49E26896";
  defparam rom_dat0_2_0_2.INITVAL_20 = "0x1F894230A207CCE1E8B8094211FC3A190E61E41000027254E51E45D27C951645617876158661E4AA";
  defparam rom_dat0_2_0_2.INITVAL_21 = "0x248EA26C6A288FE184FE0F8AA308A73E8332DC983B8EE3A88B2B4E3234E23744E3C0FA128171E0B4";
  defparam rom_dat0_2_0_2.INITVAL_22 = "0x180BA3842F02CCE3C8BF2ECA63C0AB32C8A2A0882BCEE3E8EB2E8183B06A2A8C33203A2E8092E8BE";
  defparam rom_dat0_2_0_2.INITVAL_23 = "0x2B8BE2E0BC2F0BF3E83B3CCAB3C0EF2ACF33C8673E8EB2E83F3C8EF278AA0AC483A8CE0F8AA3308B";
  defparam rom_dat0_2_0_2.INITVAL_24 = "0x2A02A2E43A3A4BA2E02B2A43A3A4BA2E82B2BC0A2F0AA278AE2D8BA2A0EE2E0AA2E8AA2E8BF2B8BF";
  defparam rom_dat0_2_0_2.INITVAL_25 = "0x3A8A33FCA60ACEE2A8BE3A06B3EC9D2A4A7258A9074AA244A61A42A0286C2E82B0F03C0F0673A8EE";
  defparam rom_dat0_2_0_2.INITVAL_26 = "0x380B515455140000882A280DB1BCF607CE23A0BF3B8BF22C540146A04402210410A04426CFE0FCFB";
  defparam rom_dat0_2_0_2.INITVAL_27 = "0x1E8A5000000000000000000000900005000050151A8AA2082104410000031CC320886A2A8A82A0AA";
  defparam rom_dat0_2_0_2.INITVAL_28 = "0x1208822088274DD374DD38822088220DC771DC771208822088274DD374DD38822088220941D16451";
  defparam rom_dat0_2_0_2.INITVAL_29 = "0x1208822088274DD374DD38822088220DC771DC771208822088274DD374DD38822088220DC771DC77";
  defparam rom_dat0_2_0_2.INITVAL_2A = "0x318D32E42C1B07904C86318D32E42C1E42C118D324C863B0790E42C118D324C863B0790DC771DC77";
  defparam rom_dat0_2_0_2.INITVAL_2B = "0x1B07904C86318D32E42C1B07904C8634C863B0790E42C118D324C863B0790E42C118D32B07904C86";
  defparam rom_dat0_2_0_2.INITVAL_2C = "0x0E81124C9324C91140820ACFA2F8AB3ECA23A8BA08892128C22283A3ECEA0ACEA2A8A8218D32E42C";
  defparam rom_dat0_2_0_2.INITVAL_2D = "0x03CFA2A8A813000000000000000000000000000000000000170082A0EC100E8100EC120A02B00C10";
  defparam rom_dat0_2_0_2.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000008C80000000000";
  defparam rom_dat0_2_0_2.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_2.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_2.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_2.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_2.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_2.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_2.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_2.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_2.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_2.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_2.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_2.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_2.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_2.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_2.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_2.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_2.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_2.OUTREG = "BYPASSED";
  defparam rom_dat0_2_0_2.RESETMODE = "SYNC";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:58955.9-58964.2" *)
  SP16K rom_dat0_2_0_3 (
    .AD({ builder_array_muxed0_12_RED_VOTER_wire, builder_array_muxed0_11_RED_VOTER_wire, builder_array_muxed0_10_RED_VOTER_wire, builder_array_muxed0_9_RED_VOTER_wire, builder_array_muxed0_8_RED_VOTER_wire, builder_array_muxed0_7_RED_VOTER_wire, builder_array_muxed0_6_RED_VOTER_wire, builder_array_muxed0_5_RED_VOTER_wire, builder_array_muxed0_4_RED_VOTER_wire, N_103_0_RED_VOTER_wire, builder_array_muxed0_2_RED_VOTER_wire, builder_array_muxed0_1_RED_VOTER_wire, builder_array_muxed0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire }),
    .CE(VCC_0_RED_VOTER_wire),
    .CLK(sys_clk),
    .CS({ VCC_0_RED_VOTER_wire, VCC_0_RED_VOTER_wire, VCC_0_RED_VOTER_wire }),
    .DI({ GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire }),
    .DO({ rom_dat0_2_0_3_DO, rom_dat0[7:6] }),
    .RST(GND_0_0_RED_VOTER_wire),
    .WE(GND_0_0_RED_VOTER_wire)
  );
  defparam rom_dat0_2_0_3.DATA_WIDTH = "X2";
  defparam rom_dat0_2_0_3.GSR = "ENABLED";
  defparam rom_dat0_2_0_3.INITVAL_00 = "0x12088220862885A120A00A00000002200971040620402108810004822088220AC000000000000001";
  defparam rom_dat0_2_0_3.INITVAL_01 = "0x0008004065104A4220A01C8490648000C110400400004020810C431028B3070D111804100690A445";
  defparam rom_dat0_2_0_3.INITVAL_02 = "0x04400288B939C413785A100E92A42C1103028C0038C40128E0118A40684806CA90A4562185220CC8";
  defparam rom_dat0_2_0_3.INITVAL_03 = "0x1401C3B00C0005E02028118971D0D018828000002402C0C00000007088C00005B30C022000100863";
  defparam rom_dat0_2_0_3.INITVAL_04 = "0x048B20000000028210C138CAA0A8A22C4CC0888208092088220C4592DC0E2C4C0288A2388AF16C4D";
  defparam rom_dat0_2_0_3.INITVAL_05 = "0x0084F2009E204910580E024020C8040209C0A088130710C4A1230C62A83123C0A23081090082208A";
  defparam rom_dat0_2_0_3.INITVAL_06 = "0x0A4BA0280A0408822CAC1C0C1218900A038000200004709089208001102208CA21E0912080008005";
  defparam rom_dat0_2_0_3.INITVAL_07 = "0x0B8040882C060B00202201019008C00702C104AB08422304AB0200010492308423048B020090142C";
  defparam rom_dat0_2_0_3.INITVAL_08 = "0x02000104922E0A4060B80484122C810882C068B0080800406406061018851C82838044060B806406";
  defparam rom_dat0_2_0_3.INITVAL_09 = "0x22C080800405C09018AC218420B0182C082000411042901C8A328410182E0101A2E010220B0188C0";
  defparam rom_dat0_2_0_3.INITVAL_0A = "0x1A8C020800104421C824068B8064060B8042406238042088C12AC00208001049C2406A32064088C1";
  defparam rom_dat0_2_0_3.INITVAL_0B = "0x08C230882C208C30C0CF030C3030C30303030C311800030884068B2068412AC212406238064220B0";
  defparam rom_dat0_2_0_3.INITVAL_0C = "0x080921C0B20908822088238482B0482382A00000080200807231C0B08C1B0AC283C0CC07C0F0CC23";
  defparam rom_dat0_2_0_3.INITVAL_0D = "0x0282A0641220000100CD29838028CA0107209C330C84102004260013043100C24148B81886427813";
  defparam rom_dat0_2_0_3.INITVAL_0E = "0x1980D208B20680A2C0E10AC08000000080029C8222082090AC0088932422090282B00222C2012841";
  defparam rom_dat0_2_0_3.INITVAL_0F = "0x248BC2087A088CA248B2288293AC2C2C083088C8208EE1E08B2A8B01985932429328A02A4A20485A";
  defparam rom_dat0_2_0_3.INITVAL_10 = "0x2EC8A3249B020E93887824489288E92BC8B0A0B020C221AC862C8E42B82C240220A081388B21E0B8";
  defparam rom_dat0_2_0_3.INITVAL_11 = "0x2448A070242B09832C3206C2E088992A8981203A370862889025887388C82C083088B81E0BB2B822";
  defparam rom_dat0_2_0_3.INITVAL_12 = "0x0540A144992642C260011446602028098A6190263A820024400442400044214A412028060860B820";
  defparam rom_dat0_2_0_3.INITVAL_13 = "0x2200013C0009021040440A4830B842040081A49106869130A819071058A80504100865294390E425";
  defparam rom_dat0_2_0_3.INITVAL_14 = "0x02088288F60004A0E00B220A21202800000004F32086C1202928800290B0000020804F2900824021";
  defparam rom_dat0_2_0_3.INITVAL_15 = "0x14045010510501016014010910141101C81008412A8202080019C29218902A8880A0620000000004";
  defparam rom_dat0_2_0_3.INITVAL_16 = "0x018060C81A14000284222441924808220882BC22118301C863098A42648826419008A92488001CF4";
  defparam rom_dat0_2_0_3.INITVAL_17 = "0x0048126CC92000411860064920681A240F210011048A4224281284A268010500022844200640404C";
  defparam rom_dat0_2_0_3.INITVAL_18 = "0x0BCC1038272A0931881E00882184780241E3E09F2207E0981810C1F210A90783C270441048410413";
  defparam rom_dat0_2_0_3.INITVAL_19 = "0x1900B0B04A0880A028B120852160A02840118C2C130091240215450058021508800000100B21B001";
  defparam rom_dat0_2_0_3.INITVAL_1A = "0x200A00A8A420000088A00A88A2A88A02868268120E0CB068202A40E000E8020A0000000A0A20A020";
  defparam rom_dat0_2_0_3.INITVAL_1B = "0x080AA2082A2082A2082A28800028000043A000022982024828240A228816288120B0041000000802";
  defparam rom_dat0_2_0_3.INITVAL_1C = "0x0248828828240230C020204080804000069020861086410088144400802011400200801608002000";
  defparam rom_dat0_2_0_3.INITVAL_1D = "0x190022A885020B01A8AA2A862020C608080084981A8622606A18892090830108420C1208001040B0";
  defparam rom_dat0_2_0_3.INITVAL_1E = "0x0A80201832058F02641A2C84C260A30849008888220B038014208B830C81020A6248000000000046";
  defparam rom_dat0_2_0_3.INITVAL_1F = "0x00028004CA298AA390100882830CCA080C002481000B30303C2880E000B8008010000B030C130000";
  defparam rom_dat0_2_0_3.INITVAL_20 = "0x0142A0A859280A809000068BA2282506093010020A0B032032030801A8E02308B0842922433030C0";
  defparam rom_dat0_2_0_3.INITVAL_21 = "0x14445154441500005000000451445A35C2A16C0022088244E500010110F90B88900887010280304A";
  defparam rom_dat0_2_0_3.INITVAL_22 = "0x15055114101145515444144151504514405144401545414040144500144000001154551544514414";
  defparam rom_dat0_2_0_3.INITVAL_23 = "0x10044154551544411411154551504505455154550545001044010000441515444154550545405445";
  defparam rom_dat0_2_0_3.INITVAL_24 = "0x14415044151545504415144151445515455054451545115055154151505505055054550545510055";
  defparam rom_dat0_2_0_3.INITVAL_25 = "0x01440004540401405401100551440100400050000140000004100141145505055054150544514455";
  defparam rom_dat0_2_0_3.INITVAL_26 = "0x1B485154551545500005150040000510001154000540001010114100501501405040501400110000";
  defparam rom_dat0_2_0_3.INITVAL_27 = "0x11045100000000000000000000000010000100000000002CBB2CC3B0CC320A8220882E2A8AB2A49E";
  defparam rom_dat0_2_0_3.INITVAL_28 = "0x2503E2503E2046B3046B3046B3046B3ACC11ACC11ACC11ACC11F8940F8940F8940F8940145114455";
  defparam rom_dat0_2_0_3.INITVAL_29 = "0x0F8940F8940ACC11ACC11ACC11ACC11046B3046B3046B3046B3503E2503E2503E2503E2503E2503E";
  defparam rom_dat0_2_0_3.INITVAL_2A = "0x0DC771DC77174DD374DD32088220882208822088274DD374DD3DC771DC7718822088220F8940F894";
  defparam rom_dat0_2_0_3.INITVAL_2B = "0x0DC771DC77174DD374DD32088220882208822088274DD374DD3DC771DC7718822088220882208822";
  defparam rom_dat0_2_0_3.INITVAL_2C = "0x0FC3C3F8A91500114455154511541414455140540045110051010151445500044040400882208822";
  defparam rom_dat0_2_0_3.INITVAL_2D = "0x13CFA2A8AA314000040000400004000040000400004000042A0A8160F03C0A42B0581500C1705802";
  defparam rom_dat0_2_0_3.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000004CC0000010000";
  defparam rom_dat0_2_0_3.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_3.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_3.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_3.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_3.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_3.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_3.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_3.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_3.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_3.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_3.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_3.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_3.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_3.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_3.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_3.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_3.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_3.OUTREG = "BYPASSED";
  defparam rom_dat0_2_0_3.RESETMODE = "SYNC";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:58874.9-58883.2" *)
  SP16K rom_dat0_2_0_4 (
    .AD({ builder_array_muxed0_12_RED_VOTER_wire, builder_array_muxed0_11_RED_VOTER_wire, builder_array_muxed0_10_RED_VOTER_wire, builder_array_muxed0_9_RED_VOTER_wire, builder_array_muxed0_8_RED_VOTER_wire, builder_array_muxed0_7_RED_VOTER_wire, builder_array_muxed0_6_RED_VOTER_wire, builder_array_muxed0_5_RED_VOTER_wire, builder_array_muxed0_4_RED_VOTER_wire, N_103_0_RED_VOTER_wire, builder_array_muxed0_2_RED_VOTER_wire, builder_array_muxed0_1_RED_VOTER_wire, builder_array_muxed0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire }),
    .CE(VCC_0_RED_VOTER_wire),
    .CLK(sys_clk),
    .CS({ VCC_0_RED_VOTER_wire, VCC_0_RED_VOTER_wire, VCC_0_RED_VOTER_wire }),
    .DI({ GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire }),
    .DO({ rom_dat0_2_0_4_DO, rom_dat0[9:8] }),
    .RST(GND_0_0_RED_VOTER_wire),
    .WE(GND_0_0_RED_VOTER_wire)
  );
  defparam rom_dat0_2_0_4.DATA_WIDTH = "X2";
  defparam rom_dat0_2_0_4.GSR = "ENABLED";
  defparam rom_dat0_2_0_4.INITVAL_00 = "0x0540F294032FC8002CBB320880A8223D4C005041150920A4541541F280FA17C81088220882200000";
  defparam rom_dat0_2_0_4.INITVAL_01 = "0x220020100A04002140D108020030E00086610822194A2078EA0104228C00220AA0844A00080200A8";
  defparam rom_dat0_2_0_4.INITVAL_02 = "0x2A088320C00C80A00C80288803F0022A8800C00020000000B202008000AC208C0000280000800090";
  defparam rom_dat0_2_0_4.INITVAL_03 = "0x220410C822020033285200CE0000052F890230EC394311208A02450168000000C050290640408C2C";
  defparam rom_dat0_2_0_4.INITVAL_04 = "0x00C8D208222541234414010AB16CBA3101111C671E4C73A4401182C3005B018043CCDF0ECD222032";
  defparam rom_dat0_2_0_4.INITVAL_05 = "0x1CC12114A2340C41ACC30F0540146114042150C5084042104408813370860A097084500C4503E850";
  defparam rom_dat0_2_0_4.INITVAL_06 = "0x158CE3B4BB11CA5000C128C18188C33648022095214000C4000202100494010D7214C60246200810";
  defparam rom_dat0_2_0_4.INITVAL_07 = "0x1C49125001130C0218582444C1502510451050DC25040058CC29841050C305410050CC2185C14041";
  defparam rom_dat0_2_0_4.INITVAL_08 = "0x21851050C3228B113CC613C1437064150011B4C2264201143113030388C0014AF06431138C613053";
  defparam rom_dat0_2_0_4.INITVAL_09 = "0x37086120111006416C7214C140044D32064204140509C148070583814C712444C31846140050CC0A";
  defparam rom_dat0_2_0_4.INITVAL_0A = "0x2DC0A190810500F014A11B8C6130531C4993143B06419100143700A19081050C1114B70943110014";
  defparam rom_dat0_2_0_4.INITVAL_0B = "0x15054168511941411410144141441414445050400E08906851134C9134163709431437064B114005";
  defparam rom_dat0_2_0_4.INITVAL_0C = "0x164EF018491C4503E85006CBC3C48D34C212E0882C0A202405060941604C15051014111005011054";
  defparam rom_dat0_2_0_4.INITVAL_0D = "0x154430B8E41282104CB8164CB27C2B308052C06E014BE3D0F2330140D04437079210CF0BC3B30C44";
  defparam rom_dat0_2_0_4.INITVAL_0E = "0x0CC7201CC63BC53310063E0642882A08C913C0CF338CF2C0F218C5C05054000BC3C8631705903400";
  defparam rom_dat0_2_0_4.INITVAL_0F = "0x100E1194012BC1F00CC03CC5C230511185805C160901B018BE3ECEF0EC8C0C0C205C8C330FB22CAE";
  defparam rom_dat0_2_0_4.INITVAL_10 = "0x3B8EF0504C1581C09401100CE2CC303C014064C616059038D3314323C4733147E240102ECC50BCC1";
  defparam rom_dat0_2_0_4.INITVAL_11 = "0x330CC10C523C44601045030F2148CE330C20B8AA004620A88A28CB00140531858164210246C2C050";
  defparam rom_dat0_2_0_4.INITVAL_12 = "0x1004B200E83A0F223C50008323F42B2CCB208CB20A8F11C0143107114C99360000BC3F22CCB3C475";
  defparam rom_dat0_2_0_4.INITVAL_13 = "0x37821040481C40413C111E0B81CC101008D2F0C63B43C088F72C42C188EF2041013C382C0882B002";
  defparam rom_dat0_2_0_4.INITVAL_14 = "0x140FA1008B040A7024841682C2C49E0A08209084310120440230CA11C40A028852E4181C45000442";
  defparam rom_dat0_2_0_4.INITVAL_15 = "0x2003000C023804408CC1044CC3C000000F03FCBE3ACEB01485060543CCEC244ED030BB2208A08811";
  defparam rom_dat0_2_0_4.INITVAL_16 = "0x1C4D0328A20B0F1170D4030CA214503E85006016064012140C144800A0033A046030022A8B402080";
  defparam rom_dat0_2_0_4.INITVAL_17 = "0x3707421014200F32C823328841100C1BC850C406330031F0C001400020F022CBF14033200211143B";
  defparam rom_dat0_2_0_4.INITVAL_18 = "0x1082414CF037CC60588938C7E2B027238C3214401702114441070C8144400040110C002F0020506E";
  defparam rom_dat0_2_0_4.INITVAL_19 = "0x084EC104192501203CC638C0F030C12A0220D0410048C2F023080020880B004682A081044050C084";
  defparam rom_dat0_2_0_4.INITVAL_1A = "0x3FCBF3E8A125CFD3A8B73E89A3FCDF3FC30330272341010C043008204C8C2DCAC30C443BCCE0C4F3";
  defparam rom_dat0_2_0_4.INITVAL_1B = "0x2F8FF3ECFF3BCBF3ECFF3ECAA2BCAA2E06F3FCDE184E72A80F21CFB3DC83258C5108D30745626CFE";
  defparam rom_dat0_2_0_4.INITVAL_1C = "0x158EC3EC2F314401245821056264162589C158E3054B1054DF220380B837080E02E0DF03CEA2F8EA";
  defparam rom_dat0_2_0_4.INITVAL_1D = "0x0CC2B3FCE81402D0547F3F4AB368023C422090CD0A8322342A0C88402CF408CFB3702F0283411409";
  defparam rom_dat0_2_0_4.INITVAL_1E = "0x150212484528C062300511411130D8250C4150FA140050646904480050562246B3A0C82288808413";
  defparam rom_dat0_2_0_4.INITVAL_1F = "0x224502108F3CCF7044451A4400501A254061F05818CC0144412A45219CEE08CDA0CC8C1441606824";
  defparam rom_dat0_2_0_4.INITVAL_20 = "0x2E0BF0FC0E3AC9C3C01133CEC1A43033CC41445E24005058452446623C1928468170F41784414408";
  defparam rom_dat0_2_0_4.INITVAL_21 = "0x1C03E0E0A72B45539C55004800000F3C8EF03CB33B0EC3001003CE30C06435CE815CF01C87F3E8BB";
  defparam rom_dat0_2_0_4.INITVAL_22 = "0x000FC19412230A20A885200250A0442304111C00380071705C040080302C00001164E93204501857";
  defparam rom_dat0_2_0_4.INITVAL_23 = "0x000A73248A22839154160A0800A0BA0D42A0A4CD2C090000C8018000ECB123084008400706908C8D";
  defparam rom_dat0_2_0_4.INITVAL_24 = "0x11415354170882535C373941409404258D520881028AD010012C8142241A050BA0144901466000A6";
  defparam rom_dat0_2_0_4.INITVAL_25 = "0x1D002280820900B034442C0150143430CCD07CC30F0FC0CC0330C3233045048C10280A0283928C11";
  defparam rom_dat0_2_0_4.INITVAL_26 = "0x040090E483260390C8133B431354503D45117C55138D5134EC14CE213C11144CD0440C3545434456";
  defparam rom_dat0_2_0_4.INITVAL_27 = "0x3C86300000000000000000000008AA20455100000000000411044110441104411044162A8A92A4BA";
  defparam rom_dat0_2_0_4.INITVAL_28 = "0x25455100000FCFF3A8AA25455100000FCFF3A8AA25455100000FCFF3A8AA25455100000FCFF3FCFF";
  defparam rom_dat0_2_0_4.INITVAL_29 = "0x30000054551A8AA2FCFF30000054551A8AA2FCFF30000054551A8AA2FCFF30000054551FCFF3A8AA";
  defparam rom_dat0_2_0_4.INITVAL_2A = "0x10441104411044110441104411044115014050140501405014050140501405014050140A8AA2FCFF";
  defparam rom_dat0_2_0_4.INITVAL_2B = "0x2F8BE2F8BE2F8BE2F8BE2F8BE2F8BE2ACEB3ACEB3ACEB3ACEB3ACEB3ACEB3ACEB3ACEB3044110441";
  defparam rom_dat0_2_0_4.INITVAL_2C = "0x05016000000000228CDF1B8923A82C3003604C80080911045100007108FD00078080800F8BE2F8BE";
  defparam rom_dat0_2_0_4.INITVAL_2D = "0x13CF00000020800000000000000000000000000000000000290A42A05C1705C1405C14054280A42A";
  defparam rom_dat0_2_0_4.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000060000010000";
  defparam rom_dat0_2_0_4.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_4.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_4.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_4.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_4.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_4.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_4.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_4.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_4.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_4.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_4.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_4.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_4.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_4.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_4.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_4.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_4.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_4.OUTREG = "BYPASSED";
  defparam rom_dat0_2_0_4.RESETMODE = "SYNC";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:58793.9-58802.2" *)
  SP16K rom_dat0_2_0_5 (
    .AD({ builder_array_muxed0_12_RED_VOTER_wire, builder_array_muxed0_11_RED_VOTER_wire, builder_array_muxed0_10_RED_VOTER_wire, builder_array_muxed0_9_RED_VOTER_wire, builder_array_muxed0_8_RED_VOTER_wire, builder_array_muxed0_7_RED_VOTER_wire, builder_array_muxed0_6_RED_VOTER_wire, builder_array_muxed0_5_RED_VOTER_wire, builder_array_muxed0_4_RED_VOTER_wire, N_103_0_RED_VOTER_wire, builder_array_muxed0_2_RED_VOTER_wire, builder_array_muxed0_1_RED_VOTER_wire, builder_array_muxed0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire }),
    .CE(VCC_0_RED_VOTER_wire),
    .CLK(sys_clk),
    .CS({ VCC_0_RED_VOTER_wire, VCC_0_RED_VOTER_wire, VCC_0_RED_VOTER_wire }),
    .DI({ GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire }),
    .DO({ rom_dat0_2_0_5_DO, rom_dat0[11:10] }),
    .RST(GND_0_0_RED_VOTER_wire),
    .WE(GND_0_0_RED_VOTER_wire)
  );
  defparam rom_dat0_2_0_5.DATA_WIDTH = "X2";
  defparam rom_dat0_2_0_5.GSR = "ENABLED";
  defparam rom_dat0_2_0_5.INITVAL_00 = "0x03CFA2A859154FA288BB07016018F43C4400504915051354541400F3E85514000014AF014AF00000";
  defparam rom_dat0_2_0_5.INITVAL_01 = "0x140A8210AD048AB3FCA20A8381C03A16CB821037268FD18C0E1D05B3E095334DF3C897028E93A8B8";
  defparam rom_dat0_2_0_5.INITVAL_02 = "0x15050088181080C1C07A0CC68000AF1ECDA220AA2A01A028C3018AD1E830320280A47A208462A01A";
  defparam rom_dat0_2_0_5.INITVAL_03 = "0x214411645110492268A63747030405368A51504519851130162F41015400000040505D1647010417";
  defparam rom_dat0_2_0_5.INITVAL_04 = "0x1388A0D45A358141041405055154551101115455154422A894110441005911815154552745131013";
  defparam rom_dat0_2_0_5.INITVAL_05 = "0x144161147D140441744D05014114501444115454084042109A3881115C8639095384551405F2A8A4";
  defparam rom_dat0_2_0_5.INITVAL_06 = "0x1546D15455008AA1485119415144452A887304A9190001405315444040A91105531445168B5258C0";
  defparam rom_dat0_2_0_5.INITVAL_07 = "0x244502A4411944C1546D0046405014104510585415014050543945C0584105404050543D41416001";
  defparam rom_dat0_2_0_5.INITVAL_08 = "0x1546005841194511944519416190540A441158413544501491110101844E19455054D11984511059";
  defparam rom_dat0_2_0_5.INITVAL_09 = "0x190E5164C1180541645116409104561385527016050A414859054D4164911446511442294052543C";
  defparam rom_dat0_2_0_5.INITVAL_0A = "0x16407154140580501451194451905924452114990540A25016190C71541405841114950549025015";
  defparam rom_dat0_2_0_5.INITVAL_0B = "0x150541545115414114101441414414144450504407014054611D4451D4161505611499054D029405";
  defparam rom_dat0_2_0_5.INITVAL_0C = "0x1544511445140FF2A8A5064541447A2B4262B01416CE614005050541507416056014111805011054";
  defparam rom_dat0_2_0_5.INITVAL_0D = "0x058911585925C04084161645519495108051407B1145B1BC621D0250B4471E06119C651541112448";
  defparam rom_dat0_2_0_5.INITVAL_0E = "0x05452114462D455114151505839C0B1742814C451DC45040511445405029104541445115055354C4";
  defparam rom_dat0_2_0_5.INITVAL_0F = "0x1146115405154151C441144541505111454154151D41D0145515445164B4390560589B15055154B5";
  defparam rom_dat0_2_0_5.INITVAL_10 = "0x19075050841541409405100572541416054164451505525C5111413144551086A294200744501445";
  defparam rom_dat0_2_0_5.INITVAL_11 = "0x1D0452085314445210450949215875154471D4452047517467194520541511454154450245524455";
  defparam rom_dat0_2_0_5.INITVAL_12 = "0x14C55320641505B1145A1E0990F4B514451164DD15459160141D0501449D120500D4D50544D14455";
  defparam rom_dat0_2_0_5.INITVAL_13 = "0x1905006055040441141105454144041D0541504515434154D534434154551C410154D41404415026";
  defparam rom_dat0_2_0_5.INITVAL_14 = "0x27CAA250171946A31454154E9198A41646F000C41545101446154EC1400739C55060241409501497";
  defparam rom_dat0_2_0_5.INITVAL_15 = "0x1145C154C718489294A218C6917044148A41545601CFC2945B0405C2A8692D8470DC593046B014C0";
  defparam rom_dat0_2_0_5.INITVAL_16 = "0x144931145D2945515C951944510C7F2A8A50F05509C5E3141815477310F61D0CD364761545D16CF1";
  defparam rom_dat0_2_0_5.INITVAL_17 = "0x250641341415451164151D4492F4653544527C6F11459150552D43519C5415456154D91541111496";
  defparam rom_dat0_2_0_5.INITVAL_18 = "0x00C101745235445154450404524C1410C05334481543314C551584C154D411CE1104331507105055";
  defparam rom_dat0_2_0_5.INITVAL_19 = "0x37454144092A452154441049501469150413505104406050412C48404841238A92C46C0140524450";
  defparam rom_dat0_2_0_5.INITVAL_1A = "0x1545515451154551545515455154551541A118A515414124A61A002164A515455154661546516459";
  defparam rom_dat0_2_0_5.INITVAL_1B = "0x1445511415144551141515455154551507515455174551D4A511455154451544110C410545515455";
  defparam rom_dat0_2_0_5.INITVAL_1C = "0x05444144151044411455140551541515414154510549105455010550505504454144550105511415";
  defparam rom_dat0_2_0_5.INITVAL_1D = "0x0441515458094051545515495154011585014C45154111145504441134540545D15005178D010405";
  defparam rom_dat0_2_0_5.INITVAL_1E = "0x1646E108851B4051D0DE1142119064150831FCAA29405054473B88C050561E8AE1A49C058C631011";
  defparam rom_dat0_2_0_5.INITVAL_1F = "0x1B4552C05514459044411A89105015154151549B2544014441154521545510464144141441508CA5";
  defparam rom_dat0_2_0_5.INITVAL_20 = "0x1505505415154561481D0D46615493194481409A29405054451445535415184581649929C8414401";
  defparam rom_dat0_2_0_5.INITVAL_21 = "0x0CCCC000300FCFF268FF0E0041801514C55014991586710010214592487515454154531485517455";
  defparam rom_dat0_2_0_5.INITVAL_22 = "0x0303F1541A0103003CC4000F503074240C71CCB0000782449616C002800000083268590EC0604064";
  defparam rom_dat0_2_0_5.INITVAL_23 = "0x120243080300C400341003005030E33D40F03C1111010000000B8000EC301C004100910045001C00";
  defparam rom_dat0_2_0_5.INITVAL_24 = "0x1C825044140000504C340341403405390F5140CE10CFA1DC41330D43489C350FD0AC5D0AC6612026";
  defparam rom_dat0_2_0_5.INITVAL_25 = "0x144B020CF0030102D841020211282F3FCCB3BCC20B0FC088033083133456284DD00C0300C2033C23";
  defparam rom_dat0_2_0_5.INITVAL_26 = "0x00005100640184000C333F4242FCF33BCF137CFF320BF3288828CA4208221848E0C80807CFC2CCFE";
  defparam rom_dat0_2_0_5.INITVAL_27 = "0x294B3000000000000000000000000000000004500800800C330CC330CC330CC330CC333FCF00F0FF";
  defparam rom_dat0_2_0_5.INITVAL_28 = "0x3FCFF3FCFF3A8AA2A8AA2A8AA2A8AA25455154551545515455100000000000000000000A8AA2A8AA";
  defparam rom_dat0_2_0_5.INITVAL_29 = "0x3FCFF3FCFF3A8AA2A8AA2A8AA2A8AA25455154551545515455100000000000000000000FCFF3FCFF";
  defparam rom_dat0_2_0_5.INITVAL_2A = "0x0FCEA254400FCEA254400FCEA254400FCEA254400FCEA254400FCEA254400FCEA254400FCFF3FCFF";
  defparam rom_dat0_2_0_5.INITVAL_2B = "0x0FCEA254400FCEA254400FCEA254400FCEA254400FCEA254400FCEA254400FCEA254400FCEA25440";
  defparam rom_dat0_2_0_5.INITVAL_2C = "0x05C1700000000000081C1B8023802C30046000840CCD3000500101D2C0010084333C3C3FCEA25440";
  defparam rom_dat0_2_0_5.INITVAL_2D = "0x23CF51545531400000000000000000000000000000000000290A4290AC280AC280A0290A01705C17";
  defparam rom_dat0_2_0_5.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000020000";
  defparam rom_dat0_2_0_5.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_5.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_5.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_5.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_5.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_5.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_5.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_5.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_5.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_5.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_5.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_5.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_5.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_5.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_5.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_5.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_5.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_5.OUTREG = "BYPASSED";
  defparam rom_dat0_2_0_5.RESETMODE = "SYNC";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:58712.9-58721.2" *)
  SP16K rom_dat0_2_0_6 (
    .AD({ builder_array_muxed0_12_RED_VOTER_wire, builder_array_muxed0_11_RED_VOTER_wire, builder_array_muxed0_10_RED_VOTER_wire, builder_array_muxed0_9_RED_VOTER_wire, builder_array_muxed0_8_RED_VOTER_wire, builder_array_muxed0_7_RED_VOTER_wire, builder_array_muxed0_6_RED_VOTER_wire, builder_array_muxed0_5_RED_VOTER_wire, builder_array_muxed0_4_RED_VOTER_wire, N_103_0_RED_VOTER_wire, builder_array_muxed0_2_RED_VOTER_wire, builder_array_muxed0_1_RED_VOTER_wire, builder_array_muxed0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire }),
    .CE(VCC_0_RED_VOTER_wire),
    .CLK(sys_clk),
    .CS({ VCC_0_RED_VOTER_wire, VCC_0_RED_VOTER_wire, VCC_0_RED_VOTER_wire }),
    .DI({ GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire }),
    .DO({ rom_dat0_2_0_6_DO, rom_dat0[13:12] }),
    .RST(GND_0_0_RED_VOTER_wire),
    .WE(GND_0_0_RED_VOTER_wire)
  );
  defparam rom_dat0_2_0_6.DATA_WIDTH = "X2";
  defparam rom_dat0_2_0_6.GSR = "ENABLED";
  defparam rom_dat0_2_0_6.INITVAL_00 = "0x028AA2A8A40481038000008AA2A8A80480111C2000C0A020010000A2A8AA2A8A02A8AA2A8AA00000";
  defparam rom_dat0_2_0_6.INITVAL_01 = "0x2A8060C8A13240E00008340C326081284982E880088122086320C11040810004200000388360C808";
  defparam rom_dat0_2_0_6.INITVAL_02 = "0x22CAA0243B1F4E13A0803A0B134C020A08102C21020E2388483BC3F000E2034D3224280B07821002";
  defparam rom_dat0_2_0_6.INITVAL_03 = "0x0EC3C1880E2A84C00080110030F0C0180082882A240080A8AA2A003028D0004D3208A8020202A0C0";
  defparam rom_dat0_2_0_6.INITVAL_04 = "0x200102A8AA200A22304330C92008500CCCA10802140022A8AA0C4030C4040C091258401000D0CCCD";
  defparam rom_dat0_2_0_6.INITVAL_05 = "0x0000408400000300402420402240040281A00828310D304C010104F0001101400010010100A2A8AA";
  defparam rom_dat0_2_0_6.INITVAL_06 = "0x0041008081008AA2A4040404129880000922A8882801C080A9028A8300AA2A0821A0810002A2A883";
  defparam rom_dat0_2_0_6.INITVAL_07 = "0x090202A8A40009A2808821001008600D008300090202A1000928088100391000A100092802100024";
  defparam rom_dat0_2_0_6.INITVAL_08 = "0x28088100382004C00090200C0024080A8A40009A208220400C0C8C703004000001084C0009020C00";
  defparam rom_dat0_2_0_6.INITVAL_09 = "0x024A02208413C03040240800A29000268082204431C03044001002B000240B000240822A8900086A";
  defparam rom_dat0_2_0_6.INITVAL_0A = "0x0086A02088110203800C10C9020C10390200C0021080A2A840024AA02088110380C002108002A840";
  defparam rom_dat0_2_0_6.INITVAL_0B = "0x0140500054014450444D05045050450505111422128A82000C10080240C4020080C402008002A890";
  defparam rom_dat0_2_0_6.INITVAL_0C = "0x084901009A080AA2A8AA210420104029000028AA22882220C001C230000001005004441241D04405";
  defparam rom_dat0_2_0_6.INITVAL_0D = "0x028AA2C4900A8A8300440000000400038C007009000600000E04801104100000210010000040D030";
  defparam rom_dat0_2_0_6.INITVAL_0E = "0x000C4030080303012009330A2208AA2A8A82840008820238200801B0202A290AA080200640030820";
  defparam rom_dat0_2_0_6.INITVAL_0F = "0x22080014F000002040B008008100202001820840088243C000300450000310C05120001008118003";
  defparam rom_dat0_2_0_6.INITVAL_10 = "0x224A202C38040EB008C02E8AA0A8E809008200800640000CAC2082E0880E2082A2A8831A08238880";
  defparam rom_dat0_2_0_6.INITVAL_11 = "0x200002C02E080B03A0002A8200A0892040A188080C0A6228120180D00820200180003A300BA08028";
  defparam rom_dat0_2_0_6.INITVAL_12 = "0x004201CC2308C040C000180483001001C04100041C00010032000003200001C0E388882682008010";
  defparam rom_dat0_2_0_6.INITVAL_13 = "0x308A83C0CA080A00700C080013080A304A40CC01000C011000000D00500000000080C320C0304080";
  defparam rom_dat0_2_0_6.INITVAL_14 = "0x228AA2A8D8030C000030000130000E2A8AA28C4120062020A1300A82808A2A8282A0C40808A24000";
  defparam rom_dat0_2_0_6.INITVAL_15 = "0x1E83728C7937832048DC2300E32CBB28408218B20000000000300010100200021244382A8AA2A880";
  defparam rom_dat0_2_0_6.INITVAL_16 = "0x2F4202C08211C780342B030D00082A2A8AA2100001020000C3000E424C0024C010C0E10CC211D00E";
  defparam rom_dat0_2_0_6.INITVAL_17 = "0x0BC0B0C0030582D010C81400004000074000C01037474000D7134453305D244DC2B03305C4D1D430";
  defparam rom_dat0_2_0_6.INITVAL_18 = "0x0906001001000011000400000200100003000034000D00300C030F4010370C0000CCCC1DC0E35CCC";
  defparam rom_dat0_2_0_6.INITVAL_19 = "0x20000000082A889250000AC1C1245400C2830000340AC1CC6B044422006B050002A8A8020B0110A0";
  defparam rom_dat0_2_0_6.INITVAL_1A = "0x17C1735C500C0C504CC401CD01F0101F0D50C010080000C49500CA22544103C340C0A51246509054";
  defparam rom_dat0_2_0_6.INITVAL_1B = "0x0108701087010870108700487004870001121C0004001380001C05411400004022B80C00C303147C";
  defparam rom_dat0_2_0_6.INITVAL_1C = "0x080AA068A0380AB0A08008C21014C9014D20943C22080030310E06A208A0384AA028820C48701087";
  defparam rom_dat0_2_0_6.INITVAL_1D = "0x33085130D00A8900E05433400004D40102A24830084C81C021320422901B1901403C50128B0000A8";
  defparam rom_dat0_2_0_6.INITVAL_1E = "0x200282303001C40220042C0CC0780B20C020A8AA2A8A0310860003120C09180062100A2A8AA2A00C";
  defparam rom_dat0_2_0_6.INITVAL_1F = "0x2A08028CCA2B813330A00A8AA22CC30CCA2224042A0B6020BC0CC3A0A0B22A029220AA0B08822882";
  defparam rom_dat0_2_0_6.INITVAL_20 = "0x32CB220808220220B80A2309802081378B20808A2A8A2204A01A019000C00300300C03004320B0AA";
  defparam rom_dat0_2_0_6.INITVAL_21 = "0x288AB238EB3A8FF1A4FE0B8FE3C0CF284880688A288220E0612000A19C880EC20328010883000802";
  defparam rom_dat0_2_0_6.INITVAL_22 = "0x2A0962E82F128E32ECAA3382B2E0F83B88A2A0403ACEA2B4AB2A8A03B888238F2380F21088E0ECAA";
  defparam rom_dat0_2_0_6.INITVAL_23 = "0x3BCCA2B8EE3B8EE3A82B2E0EF2E09F3A8BA2E4FA3E8E33F87F3C0FF208EA3B8C83ACA20B8AE278CA";
  defparam rom_dat0_2_0_6.INITVAL_24 = "0x2A82A3A82A2EC3A3A82B2E8283E83B2ECAA3AC8B2B8E72ECAE3FCE82F0AF3A0AA2A8BA2A88B3BCCB";
  defparam rom_dat0_2_0_6.INITVAL_25 = "0x2EC433E8A808CFC2AC3F320FA2B89B154A63A8690685A244A91A42A22CBA2A8BA0B82E0B81F3F82A";
  defparam rom_dat0_2_0_6.INITVAL_26 = "0x2A8AF3FC00000000C8222A89F1BCFE27CE32A8BF3907F200542304A0D42A23440000D43ACFE1ACF8";
  defparam rom_dat0_2_0_6.INITVAL_27 = "0x2B8A000000000000000000000010000500005005128AA28000000000000000000000091545A25855";
  defparam rom_dat0_2_0_6.INITVAL_28 = "0x34C9324C932B06C1B06C1E4390E439018C6318C634C9324C932B06C1B06C1E4390E4390A8AA2A8AA";
  defparam rom_dat0_2_0_6.INITVAL_29 = "0x218C6318C63E4390E4390B06C1B06C14C9324C93218C6318C63E4390E4390B06C1B06C118C6318C6";
  defparam rom_dat0_2_0_6.INITVAL_2A = "0x3C4B12C4B12384E1384E16C1B06C1B090E4390E43C4B12C4B12384E1384E16C1B06C1B04C9324C93";
  defparam rom_dat0_2_0_6.INITVAL_2B = "0x3C4B12C4B12384E1384E16C1B06C1B090E4390E43C4B12C4B12384E1384E16C1B06C1B090E4390E4";
  defparam rom_dat0_2_0_6.INITVAL_2C = "0x000000000000000000E322CE82FC8A2A8FB3ACFE088A2238A22383A28CEE08CB222828290E4390E4";
  defparam rom_dat0_2_0_6.INITVAL_2D = "0x03CF0000000280000000000000000000000000000000000001004000000100001004010040000000";
  defparam rom_dat0_2_0_6.INITVAL_2E = "0x000000000000000000000000000000000000000000000000000000000000000000040F0000000000";
  defparam rom_dat0_2_0_6.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_6.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_6.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_6.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_6.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_6.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_6.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_6.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_6.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_6.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_6.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_6.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_6.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_6.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_6.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_6.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_6.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_6.OUTREG = "BYPASSED";
  defparam rom_dat0_2_0_6.RESETMODE = "SYNC";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:58631.9-58640.2" *)
  SP16K rom_dat0_2_0_7 (
    .AD({ builder_array_muxed0_12_RED_VOTER_wire, builder_array_muxed0_11_RED_VOTER_wire, builder_array_muxed0_10_RED_VOTER_wire, builder_array_muxed0_9_RED_VOTER_wire, builder_array_muxed0_8_RED_VOTER_wire, builder_array_muxed0_7_RED_VOTER_wire, builder_array_muxed0_6_RED_VOTER_wire, builder_array_muxed0_5_RED_VOTER_wire, builder_array_muxed0_4_RED_VOTER_wire, N_103_0_RED_VOTER_wire, builder_array_muxed0_2_RED_VOTER_wire, builder_array_muxed0_1_RED_VOTER_wire, builder_array_muxed0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire }),
    .CE(VCC_0_RED_VOTER_wire),
    .CLK(sys_clk),
    .CS({ VCC_0_RED_VOTER_wire, VCC_0_RED_VOTER_wire, VCC_0_RED_VOTER_wire }),
    .DI({ GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire }),
    .DO({ rom_dat0_2_0_7_DO, rom_dat0[15:14] }),
    .RST(GND_0_0_RED_VOTER_wire),
    .WE(GND_0_0_RED_VOTER_wire)
  );
  defparam rom_dat0_2_0_7.DATA_WIDTH = "X2";
  defparam rom_dat0_2_0_7.GSR = "ENABLED";
  defparam rom_dat0_2_0_7.INITVAL_00 = "0x20000000042A8AE1A02000000000000002000C0200C0001800000000000000004000000000000000";
  defparam rom_dat0_2_0_7.INITVAL_01 = "0x0002A2C8EA328E600008388CB2880A080000E888000822282128C232A0A2020A120008388B10E48E";
  defparam rom_dat0_2_0_7.INITVAL_02 = "0x22CAA0A8BB2F8E2370EE1A07A32C200103802408028E23A8A839CBD2B8620B8CB2A8B72B0B208802";
  defparam rom_dat0_2_0_7.INITVAL_03 = "0x0E03020000000000000202C0003001280002882201890100000001308010000600100220402000E0";
  defparam rom_dat0_2_0_7.INITVAL_04 = "0x0544400000010281300708CE701CA110C0301C070946000000008A700018200121ECA52A8130C0C0";
  defparam rom_dat0_2_0_7.INITVAL_05 = "0x000AA3002B2A0B20A42A2000400040040000A804308CB00CA00000F2C0080002C100932001000000";
  defparam rom_dat0_2_0_7.INITVAL_06 = "0x1984A028200800000820000282A80019040000140109E0200020440320000088802000208000500B";
  defparam rom_dat0_2_0_7.INITVAL_07 = "0x00028000001B0000008200070010001C042318C000800018C00002001C3801080018C00002805800";
  defparam rom_dat0_2_0_7.INITVAL_08 = "0x0002001C322088C1B000080C630002000001B00000008004CC1E8EB038A0080000088C1B00028C1B";
  defparam rom_dat0_2_0_7.INITVAL_09 = "0x300000080017C0306C00020800006C000000800531C43068880082306C000306C00020000012C000";
  defparam rom_dat0_2_0_7.INITVAL_0A = "0x2C00000020014A03200C1B00008C1B000080C4B00008000006300000002001C300C4B00008800006";
  defparam rom_dat0_2_0_7.INITVAL_0B = "0x0100408050214040040C04004040040404101005200003080C1B0000C0C6300020C4B00008800001";
  defparam rom_dat0_2_0_7.INITVAL_0C = "0x2800C0000202000000000283024008168A82000008008000C808C030002401085004001301C00004";
  defparam rom_dat0_2_0_7.INITVAL_0D = "0x020010E020080003080A32426028100B8C807084020101140E0B0200040010092000282C0082C830";
  defparam rom_dat0_2_0_7.INITVAL_0E = "0x00048298000B41210002110000800000010268AA08820238A00A01B00800000262802806002308A0";
  defparam rom_dat0_2_0_7.INITVAL_0F = "0x00020214FA000380203B020002A0000009008002220883E0023E854220E322CE80008A188A2148B1";
  defparam rom_dat0_2_0_7.INITVAL_10 = "0x0880800CF0060C3080C80CC03200C02208008000240082A40E0008C200CC0800000003208003E008";
  defparam rom_dat0_2_0_7.INITVAL_11 = "0x288600C00C20030300020CC82000220A820120283C00A008202C00E0800800090020903203320800";
  defparam rom_dat0_2_0_7.INITVAL_12 = "0x028201CC9B26C180D0810C4EE3003006C18000182F8101088E308080EC0800C9E388202E82608020";
  defparam rom_dat0_2_0_7.INITVAL_13 = "0x33000358400A00201C8C0480312080380042DCA8380EA280AB020E222CE002082080C322C2300882";
  defparam rom_dat0_2_0_7.INITVAL_14 = "0x000000006C010E0228900A8332208C0000000C60210482080230C002600000008040C62A00000422";
  defparam rom_dat0_2_0_7.INITVAL_15 = "0x0D41314434134311284C1380713C77140B4000D10000000000390282C80C00009044B10000000008";
  defparam rom_dat0_2_0_7.INITVAL_16 = "0x274A00E0210141420CAB2104008080000000102E00018108C32204A20C8820C08248C804C110500D";
  defparam rom_dat0_2_0_7.INITVAL_17 = "0x29C2B0E40B0440C000C400000028B821C420C01833CB8180F1210EE19044104462B8110440D0D012";
  defparam rom_dat0_2_0_7.INITVAL_18 = "0x00002088C82AC2008C62008801008802034120B42E0D20B82C030F4220BF2D0102CCCC07C2C34C44";
  defparam rom_dat0_2_0_7.INITVAL_19 = "0x3002820082000033680000C0C234B020C00320823C80C0ECC300800000410A088000002003000002";
  defparam rom_dat0_2_0_7.INITVAL_1A = "0x30C30368C824055088640A85829818090EC2E0000C8202CCE128C01104090A49402C501F49B07090";
  defparam rom_dat0_2_0_7.INITVAL_1B = "0x1D4AB354AB354AB354AB35C2115C21118C70844606003368001D0CE2C466204200300C2041C13C0C";
  defparam rom_dat0_2_0_7.INITVAL_1C = "0x04800240082C0430C04820C13084C50185305414310C8250912E82A208803A0AA028002F42117421";
  defparam rom_dat0_2_0_7.INITVAL_1D = "0x3B02B2F0F2000002E8BB33C2000CD2030000CC382A8EA2E0AA3A8A0020131201802C603002208030";
  defparam rom_dat0_2_0_7.INITVAL_1E = "0x10802038302A4282A8002E0CC0980302C200000000031300612003931C040602A2B800000000008E";
  defparam rom_dat0_2_0_7.INITVAL_1F = "0x0004200CC0038293B0701000031CE0084E21080C2A0370707E0081E0903A2A028220A3078C430020";
  defparam rom_dat0_2_0_7.INITVAL_20 = "0x10C380E0A2080220382023828200881983306000000313247017096228C2038032AC230003B070C0";
  defparam rom_dat0_2_0_7.INITVAL_21 = "0x1445505045150001540005454148EF020882B08A088220C8822000000C220CC22008080087800000";
  defparam rom_dat0_2_0_7.INITVAL_22 = "0x01055154101105105045100550504405005154501444515404144041101400001144011444505455";
  defparam rom_dat0_2_0_7.INITVAL_23 = "0x10045114451145105415050450505405415054551505000040050000445115044104510545505445";
  defparam rom_dat0_2_0_7.INITVAL_24 = "0x15415154150441515415154141541515455144451141511045044141545105055054550544010040";
  defparam rom_dat0_2_0_7.INITVAL_25 = "0x11450004510501505441140151141515405000410405004401104111145404455014050141404411";
  defparam rom_dat0_2_0_7.INITVAL_26 = "0x00000000551545504001150141000114001154000040001054104450141100445050141400004000";
  defparam rom_dat0_2_0_7.INITVAL_27 = "0x01411000000000000000000000000010000100000800000411044110441104411044100000000000";
  defparam rom_dat0_2_0_7.INITVAL_28 = "0x1A8BF300151A8BF300151A8BF300151FCEA254400FCEA254400FCEA254400FCEA254400000000000";
  defparam rom_dat0_2_0_7.INITVAL_29 = "0x300151A8BF300151A8BF300151A8BF354400FCEA254400FCEA254400FCEA254400FCEA2A8BF30015";
  defparam rom_dat0_2_0_7.INITVAL_2A = "0x1502B3F8811502B3F8811502B3F8811047E2ACD40047E2ACD40047E2ACD40047E2ACD4000151A8BF";
  defparam rom_dat0_2_0_7.INITVAL_2B = "0x3F8811502B3F8811502B3F8811502B3ACD40047E2ACD40047E2ACD40047E2ACD40047E2502B3F881";
  defparam rom_dat0_2_0_7.INITVAL_2C = "0x05014000000000000455100500140010054144140045111451010151145500415154541F8811502B";
  defparam rom_dat0_2_0_7.INITVAL_2D = "0x13CF5154551000000000000000000000000000000000000014050140501405014050140501405014";
  defparam rom_dat0_2_0_7.INITVAL_2E = "0x0000000000000000000000000000000000000000000000000000000000000000000C000000010000";
  defparam rom_dat0_2_0_7.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_7.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_7.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_7.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_7.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_7.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_7.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_7.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_7.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_7.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_7.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_7.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_7.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_7.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_7.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_7.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_7.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_7.OUTREG = "BYPASSED";
  defparam rom_dat0_2_0_7.RESETMODE = "SYNC";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:58550.9-58559.2" *)
  SP16K rom_dat0_2_0_8 (
    .AD({ builder_array_muxed0_12_RED_VOTER_wire, builder_array_muxed0_11_RED_VOTER_wire, builder_array_muxed0_10_RED_VOTER_wire, builder_array_muxed0_9_RED_VOTER_wire, builder_array_muxed0_8_RED_VOTER_wire, builder_array_muxed0_7_RED_VOTER_wire, builder_array_muxed0_6_RED_VOTER_wire, builder_array_muxed0_5_RED_VOTER_wire, builder_array_muxed0_4_RED_VOTER_wire, N_103_0_RED_VOTER_wire, builder_array_muxed0_2_RED_VOTER_wire, builder_array_muxed0_1_RED_VOTER_wire, builder_array_muxed0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire }),
    .CE(VCC_0_RED_VOTER_wire),
    .CLK(sys_clk),
    .CS({ VCC_0_RED_VOTER_wire, VCC_0_RED_VOTER_wire, VCC_0_RED_VOTER_wire }),
    .DI({ GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire }),
    .DO({ rom_dat0_2_0_8_DO, rom_dat0[17:16] }),
    .RST(GND_0_0_RED_VOTER_wire),
    .WE(GND_0_0_RED_VOTER_wire)
  );
  defparam rom_dat0_2_0_8.DATA_WIDTH = "X2";
  defparam rom_dat0_2_0_8.GSR = "ENABLED";
  defparam rom_dat0_2_0_8.INITVAL_00 = "0x054551545C2FC810E03300455154540146014C5504C9618411118151545515451154551545500000";
  defparam rom_dat0_2_0_8.INITVAL_01 = "0x000230CC383301B0000C300E33CC082C4992FCC0098AB32C3039C00200E002002000003CC0E00808";
  defparam rom_dat0_2_0_8.INITVAL_02 = "0x2AC000B00F330FA130812F8833CC082380803C08038F33CCFE3F008004B320C33330001C83008813";
  defparam rom_dat0_2_0_8.INITVAL_03 = "0x0C47034411154100080303C5413004300003CCFB04CC1014551544301400000300405615054150EE";
  defparam rom_dat0_2_0_8.INITVAL_04 = "0x1000215455144750701300CE701CB110C0311C671D4451545500CF710040004070FCD537C530D0D0";
  defparam rom_dat0_2_0_8.INITVAL_05 = "0x014253646B3B0F40F41F3A051110111140105411388CF23C46008031D00A0008D004430044515455";
  defparam rom_dat0_2_0_8.INITVAL_06 = "0x04C7A3F8741145515003300263EC0804401154411440F00454010153045514CE4134000245510453";
  defparam rom_dat0_2_0_8.INITVAL_07 = "0x14401154510F4451501514430144150C41034CD40405504CD41501504C3C0441504CD41507410051";
  defparam rom_dat0_2_0_8.INITVAL_08 = "0x1505504C3B2D4CD0F444000D335040154510F44514055110CD0FCFF038FF380010404D0F44404C4F";
  defparam rom_dat0_2_0_8.INITVAL_09 = "0x350540545103C5313C50100151443D114411541034C03134040808313C510743D11045154443D415";
  defparam rom_dat0_2_0_8.INITVAL_0A = "0x3D41510455040303184D0F04400C4F044000D0F50401515413350551045504C310D0F50100115413";
  defparam rom_dat0_2_0_8.INITVAL_0B = "0x1004014001100100100C10010100101040404000314553440D0F4410C0D3350100D0F50400115444";
  defparam rom_dat0_2_0_8.INITVAL_0C = "0x0C47C13447344551545513CF230C4D03CE01545511441114C105C571503410010010010704C00040";
  defparam rom_dat0_2_0_8.INITVAL_0D = "0x134541FC9E19455378F51DC2F10CB0030CD030FC010FF00C4C0C8413D44F300C41C03F2C00F3DC74";
  defparam rom_dat0_2_0_8.INITVAL_0E = "0x110C10DC440F4570140611051154551544530CFF0CC30330C11340301055140703044D0005130060";
  defparam rom_dat0_2_0_8.INITVAL_0F = "0x11041100F11487D0707F0701430010110041C400054583D44B3AC3F220E30CC21070CC0DCFB088B3";
  defparam rom_dat0_2_0_8.INITVAL_10 = "0x1DC5D01C74110D7084C01DC5405414340041C044010013F45F104DD344CD114551544335C4133440";
  defparam rom_dat0_2_0_8.INITVAL_11 = "0x0CC301CC1D34074150001D892050771F02F2F8283C072338233DC0C0041C11004004153207404014";
  defparam rom_dat0_2_0_8.INITVAL_12 = "0x084300CCFF3FC3C0FCE3180EF200230FC3C2203C2ACFD05007184110748415C0C3C0FC3B00F00074";
  defparam rom_dat0_2_0_8.INITVAL_13 = "0x3145531C55144500F40C0CC03174153D4553DCCF3D4FC3F8F5240FC3F8D4280040C0C730C3308071";
  defparam rom_dat0_2_0_8.INITVAL_14 = "0x154551542D040161241826002328591545515C711005D0505331455304451545D114C70045514017";
  defparam rom_dat0_2_0_8.INITVAL_15 = "0x3C0CF030F30F03C3C03D07C723EC3300CF33F4FE00000000003D8D71743512450100F51545515451";
  defparam rom_dat0_2_0_8.INITVAL_16 = "0x034011E061130C0104000CC3301455154551181807035184C7060100CC900CCC410013088F001CFC";
  defparam rom_dat0_2_0_8.INITVAL_17 = "0x00C030D487000CC330C30CC07100011F061310430C0043DC03170003B0C216C30000CC000CD1D4CC";
  defparam rom_dat0_2_0_8.INITVAL_18 = "0x144141FCD33744A254493B478118272D871190761E0D90740030C36100431C0181F0CC3CCCD35C73";
  defparam rom_dat0_2_0_8.INITVAL_19 = "0x22030248161544632C0A05C7E230A021C15300923845D3ECBD348831C03D39CA5154550507000454";
  defparam rom_dat0_2_0_8.INITVAL_1A = "0x3FCFF368912E0F5288670E8583DC5C3DCE83E0201C0242C82030C57144B823CF0320441F0F30E083";
  defparam rom_dat0_2_0_8.INITVAL_1B = "0x2FCEF3ECEF3BCEF3ECEF3ECAA2ECAA2F0DF3BCD611CC5108110ECDE3D4C12C0451745C0781D23CFF";
  defparam rom_dat0_2_0_8.INITVAL_1C = "0x11CD53547C2D4170D41615C45054D10545311814344C1050D11F0FF30CC43CCFF03C1D0FCAA2FCAA";
  defparam rom_dat0_2_0_8.INITVAL_1D = "0x3FC8F3F0F41547D150FF33C68010CE018551147D28CF83F4A33E0C517C1707C1F02C3C1546401075";
  defparam rom_dat0_2_0_8.INITVAL_1E = "0x05455178741F4790C0152DCDC0DC171DC050545515474314340003034C111200E29895154551540F";
  defparam rom_dat0_2_0_8.INITVAL_1F = "0x1541515C4003C35374350545534CC1110F7004023F0331343C0504F1C01F3F03D330F3130D239465";
  defparam rom_dat0_2_0_8.INITVAL_20 = "0x20CFF2EC3B380330385A23CB8100C33FC33104551547434036334A1378C0070C704C0304433130D5";
  defparam rom_dat0_2_0_8.INITVAL_21 = "0x2C47C104613F8550A45501066140FF00C8C0F0CF0CC330F0712FC0C2C41D04CA007C030C8FF32C8F";
  defparam rom_dat0_2_0_8.INITVAL_22 = "0x0D00D0400030071170CC30071270600648D06C102040B0508C0D4B4150D002000040D31408106CAF";
  defparam rom_dat0_2_0_8.INITVAL_23 = "0x1C05B2589715CB820433370550703C010DC3705E1A0500008004C0004866100401C0910C8003D4C0";
  defparam rom_dat0_2_0_8.INITVAL_24 = "0x06C340C415354140C00435C3415C14014441E4C439C423AC8515874328611502106060360401C090";
  defparam rom_dat0_2_0_8.INITVAL_25 = "0x1D010120090D4C7394A81F05C3301B3FCC6380F1030D0040C00042633088378CA09C2709C2905C3B";
  defparam rom_dat0_2_0_8.INITVAL_26 = "0x0000A2A800000000482101C0519455254520009517CD511414254451642405C4B00454324553F454";
  defparam rom_dat0_2_0_8.INITVAL_27 = "0x0201300000000000000000000008AA28455140000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_8.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_8.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_8.INITVAL_2A = "0x16C0E190F12385B0C4A43C4A43385B090F126C0E16C0E190F12385B0C4A43C4A43385B0000000000";
  defparam rom_dat0_2_0_8.INITVAL_2B = "0x16C0E190F12385B0C4A43C4A43385B090F126C0E16C0E190F12385B0C4A43C4A43385B090F126C0E";
  defparam rom_dat0_2_0_8.INITVAL_2C = "0x00000000000000000818110C0130442600410017080102005001C2000C310040111414190F126C0E";
  defparam rom_dat0_2_0_8.INITVAL_2D = "0x14CF0000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_8.INITVAL_2E = "0x0000000000000000000000000000000000000000000000000000000000000000000C003000014000";
  defparam rom_dat0_2_0_8.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_8.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_8.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_8.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_8.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_8.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_8.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_8.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_8.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_8.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_8.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_8.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_8.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_8.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_8.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_8.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_8.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_8.OUTREG = "BYPASSED";
  defparam rom_dat0_2_0_8.RESETMODE = "SYNC";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:58469.9-58478.2" *)
  SP16K rom_dat0_2_0_9 (
    .AD({ builder_array_muxed0_12_RED_VOTER_wire, builder_array_muxed0_11_RED_VOTER_wire, builder_array_muxed0_10_RED_VOTER_wire, builder_array_muxed0_9_RED_VOTER_wire, builder_array_muxed0_8_RED_VOTER_wire, builder_array_muxed0_7_RED_VOTER_wire, builder_array_muxed0_6_RED_VOTER_wire, builder_array_muxed0_5_RED_VOTER_wire, builder_array_muxed0_4_RED_VOTER_wire, N_103_0_RED_VOTER_wire, builder_array_muxed0_2_RED_VOTER_wire, builder_array_muxed0_1_RED_VOTER_wire, builder_array_muxed0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire }),
    .CE(VCC_0_RED_VOTER_wire),
    .CLK(sys_clk),
    .CS({ VCC_0_RED_VOTER_wire, VCC_0_RED_VOTER_wire, VCC_0_RED_VOTER_wire }),
    .DI({ GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire, GND_0_0_RED_VOTER_wire }),
    .DO({ rom_dat0_2_0_9_DO, rom_dat0[19:18] }),
    .RST(GND_0_0_RED_VOTER_wire),
    .WE(GND_0_0_RED_VOTER_wire)
  );
  defparam rom_dat0_2_0_9.DATA_WIDTH = "X2";
  defparam rom_dat0_2_0_9.GSR = "ENABLED";
  defparam rom_dat0_2_0_9.INITVAL_00 = "0x0000000004154692403300000000001045014C5504C5514411100000000000000000000000000000";
  defparam rom_dat0_2_0_9.INITVAL_01 = "0x2A8192C4963189D000063A8FB12086368EE3D0080EC7C0145515C221A052010A320008364A30AC8E";
  defparam rom_dat0_2_0_9.INITVAL_02 = "0x15CAA058A70B8DD240E935CA802CAE38CA6210A6214D936407368A92A4D13A08B198BE16CBA26491";
  defparam rom_dat0_2_0_9.INITVAL_03 = "0x1D470198422A850008011549413404140001445D05441000000040314000000500400114040150D5";
  defparam rom_dat0_2_0_9.INITVAL_04 = "0x0000100000044140301304C510045000C0110411140000000000453000441041115450154021C0C1";
  defparam rom_dat0_2_0_9.INITVAL_05 = "0x0141515455150740541515010014101005005400388CB22C9A0583D1600A050B6004811004000000";
  defparam rom_dat0_2_0_9.INITVAL_06 = "0x04415154100000000412150291544808800000010000D14001140003400001469118411544000003";
  defparam rom_dat0_2_0_9.INITVAL_07 = "0x1001000001054000005100410040040C411344500100004450000500443404400044500001410001";
  defparam rom_dat0_2_0_9.INITVAL_08 = "0x00090044351684D05400140D1140040000105400004440104D0D4D703455140050048D0540018C45";
  defparam rom_dat0_2_0_9.INITVAL_09 = "0x140001440103CA3114400500000415000050401034C031185809457114400B415000800000415000";
  defparam rom_dat0_2_0_9.INITVAL_0A = "0x1500001410040103288D0500014C45000140D05400400000111400001410044320D0540044000011";
  defparam rom_dat0_2_0_9.INITVAL_0B = "0x1004014001100101101C10410104101040404041100003880D05400140D1140050D0540044000004";
  defparam rom_dat0_2_0_9.INITVAL_0C = "0x14495124012800000000014561088A014651400004004000C609C070005000060010110704C11040";
  defparam rom_dat0_2_0_9.INITVAL_0D = "0x01000054551400039855154551145017CC7130A913469108CF0589329C492108724015144051D478";
  defparam rom_dat0_2_0_9.INITVAL_0E = "0x1104515400054510000111000050000080010455044101345215807000000141114856110A514454";
  defparam rom_dat0_2_0_9.INITVAL_0F = "0x00091140F6018540543511440150000144004815110443E019154151105319C65020450445504451";
  defparam rom_dat0_2_0_9.INITVAL_10 = "0x2440400CB011443080C40C409108401104004085100551540D0084C1085400080000071040035004";
  defparam rom_dat0_2_0_9.INITVAL_11 = "0x144540C80C1003510045048820009105415154141C095114111540D0400421440154503201110400";
  defparam rom_dat0_2_0_9.INITVAL_12 = "0x0C4102CC771DC940D4501C85D1001105414118141545505005144100544401C4D344541541504454";
  defparam rom_dat0_2_0_9.INITVAL_13 = "0x1100035450040000540C14411154001540415C45154D415455140D415454140040404710C1304059";
  defparam rom_dat0_2_0_9.INITVAL_14 = "0x08000000EA194D6228582A411114540000000C511504400401114001000000005000C51402005415";
  defparam rom_dat0_2_0_9.INITVAL_15 = "0x2D45B154B51B4351946E1B4E718C77148A5150190000000000398AE16424014CC030550000000000";
  defparam rom_dat0_2_0_9.INITVAL_16 = "0x174510E011354541045515462000C000000018670AC2E188F73D04D18C8418C4D3444504461178AD";
  defparam rom_dat0_2_0_9.INITVAL_17 = "0x15C170F48B0544C210C50880A25CF735462164BD15454144551D0F5150551D455154550548D1D455";
  defparam rom_dat0_2_0_9.INITVAL_18 = "0x004001545115445154450444411414114721B0B6264DB0BC1411476210D73F4D82D4FF15C7C35C55";
  defparam rom_dat0_2_0_9.INITVAL_19 = "0x1101424402000121640A0A495114A411C2A11091388A615C95144412405515455000000043010400";
  defparam rom_dat0_2_0_9.INITVAL_1A = "0x15455154511505514455054541541415CE91E050144241C8A518CA91645519455158661585906095";
  defparam rom_dat0_2_0_9.INITVAL_1B = "0x1445511455144551145515455154551505515455114451A4110D45515441140400300C0541511455";
  defparam rom_dat0_2_0_9.INITVAL_1C = "0x01455154542C4031C41510C45054D1054531141434441050511D0551044434455014140D05511455";
  defparam rom_dat0_2_0_9.INITVAL_1D = "0x3745515058000151545511494000C50144000435154D51D45535440014130141502C141402000031";
  defparam rom_dat0_2_0_9.INITVAL_1E = "0x05441038BD39859154D92E8EF164530AC003000000034364283007034C522200515450000000000D";
  defparam rom_dat0_2_0_9.INITVAL_1F = "0x0041500C95174593B4310000034CD2258D500806150331343D0A46D140251541611053134D234014";
  defparam rom_dat0_2_0_9.INITVAL_20 = "0x10C5515415140110345519454100411543310020000343543623492158D1074871844114437134C0";
  defparam rom_dat0_2_0_9.INITVAL_21 = "0x3C87D0006D378FF050FF09404240D50044405045044110D051154241641504450054010445511445";
  defparam rom_dat0_2_0_9.INITVAL_22 = "0x110910141801C4104071024551405406C03010203C40F3E88E0144825020000E00C42234CC708013";
  defparam rom_dat0_2_0_9.INITVAL_23 = "0x1380F0D404010FD34C040404A1404013011040BF0CCB020000000200CC4C0048C110510000431C08";
  defparam rom_dat0_2_0_9.INITVAL_24 = "0x0100C0100D0482C0100C0900C1901C134CC0C404310DF330373BC0C10CF103075170F4070C013800";
  defparam rom_dat0_2_0_9.INITVAL_25 = "0x04021100120304B0ACC02C0C31BC0A3FCC22C0F003CE0000C00000C33000000C0010040100304C33";
  defparam rom_dat0_2_0_9.INITVAL_26 = "0x0000F3FC000000004821170072BCFD33CF3050BF3ECBF3280007C021C0051700C084D00ACFF22CFC";
  defparam rom_dat0_2_0_9.INITVAL_27 = "0x02C10000000000000000000000000000000004500000A00000000000000000000000000000000000";
  defparam rom_dat0_2_0_9.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_9.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_9.INITVAL_2A = "0x1E047248ED048ED0E04721CB81B412348ED0E04721CB81B4123B41231CB81E047248ED0000000000";
  defparam rom_dat0_2_0_9.INITVAL_2B = "0x348ED0E0472E047248ED0B41231CB81E047248ED0B41231CB811CB81B412348ED0E0472B41231CB8";
  defparam rom_dat0_2_0_9.INITVAL_2C = "0x00000000000000000879310C4130040481C140150CC43304710143410C07004811141411CB81B412";
  defparam rom_dat0_2_0_9.INITVAL_2D = "0x20CF0000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_9.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000008000000020000";
  defparam rom_dat0_2_0_9.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_9.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_9.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_9.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_9.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_9.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_9.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_9.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_9.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_9.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_9.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_9.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_9.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_9.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_9.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_9.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_9.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
  defparam rom_dat0_2_0_9.OUTREG = "BYPASSED";
  defparam rom_dat0_2_0_9.RESETMODE = "SYNC";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55568.6-55571.2" *)
  IB serial_rx_pad (
    .I(serial_rx),
    .O(serial_rx_c)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51683.12-51689.2" *)
  OFD1P3JX serial_tx_0io_TMR_0 (
    .CK(sys_clk),
    .D(serial_tx_4_TMR_0),
    .PD(sys_rst_TMR_0),
    .Q(serial_tx_c_TMR_0),
    .SP(main_basesoc_serial_tx_rs232phytx_next_value1_1_sqmuxa_i_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51683.12-51689.2" *)
  OFD1P3JX serial_tx_0io_TMR_1 (
    .CK(sys_clk),
    .D(serial_tx_4_TMR_1),
    .PD(sys_rst_TMR_1),
    .Q(serial_tx_c_TMR_1),
    .SP(main_basesoc_serial_tx_rs232phytx_next_value1_1_sqmuxa_i_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51683.12-51689.2" *)
  OFD1P3JX serial_tx_0io_TMR_2 (
    .CK(sys_clk),
    .D(serial_tx_4_TMR_2),
    .PD(sys_rst_TMR_2),
    .Q(serial_tx_c_TMR_2),
    .SP(main_basesoc_serial_tx_rs232phytx_next_value1_1_sqmuxa_i_TMR_2)
  );
  LUT4 serial_tx_c_0_RED_VOTER (
    .A(serial_tx_c_TMR_0),
    .B(serial_tx_c_TMR_1),
    .C(serial_tx_c_TMR_2),
    .D(1'h0),
    .Z(serial_tx_c_0_RED_VOTER_wire)
  );
  defparam serial_tx_c_0_RED_VOTER.INIT = "0xFCC0";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55563.6-55566.2" *)
  OB serial_tx_pad (
    .I(serial_tx_c_0_RED_VOTER_wire),
    .O(serial_tx)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51755.11-51761.2" *)
  FD1P3IX \storage_1_dat1_reg[0]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(storage_1_TMR_0[0]),
    .Q(storage_1_dat1_TMR_0[0]),
    .SP(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51755.11-51761.2" *)
  FD1P3IX \storage_1_dat1_reg[0]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(storage_1_TMR_1[0]),
    .Q(storage_1_dat1_TMR_1[0]),
    .SP(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51755.11-51761.2" *)
  FD1P3IX \storage_1_dat1_reg[0]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(storage_1_TMR_2[0]),
    .Q(storage_1_dat1_TMR_2[0]),
    .SP(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51763.11-51769.2" *)
  FD1P3IX \storage_1_dat1_reg[1]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(storage_1_TMR_0[1]),
    .Q(storage_1_dat1_TMR_0[1]),
    .SP(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51763.11-51769.2" *)
  FD1P3IX \storage_1_dat1_reg[1]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(storage_1_TMR_1[1]),
    .Q(storage_1_dat1_TMR_1[1]),
    .SP(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51763.11-51769.2" *)
  FD1P3IX \storage_1_dat1_reg[1]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(storage_1_TMR_2[1]),
    .Q(storage_1_dat1_TMR_2[1]),
    .SP(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51771.11-51777.2" *)
  FD1P3IX \storage_1_dat1_reg[2]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(storage_1_TMR_0[2]),
    .Q(storage_1_dat1_TMR_0[2]),
    .SP(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51771.11-51777.2" *)
  FD1P3IX \storage_1_dat1_reg[2]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(storage_1_TMR_1[2]),
    .Q(storage_1_dat1_TMR_1[2]),
    .SP(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51771.11-51777.2" *)
  FD1P3IX \storage_1_dat1_reg[2]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(storage_1_TMR_2[2]),
    .Q(storage_1_dat1_TMR_2[2]),
    .SP(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51779.11-51785.2" *)
  FD1P3IX \storage_1_dat1_reg[3]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(storage_1_TMR_0[3]),
    .Q(storage_1_dat1_TMR_0[3]),
    .SP(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51779.11-51785.2" *)
  FD1P3IX \storage_1_dat1_reg[3]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(storage_1_TMR_1[3]),
    .Q(storage_1_dat1_TMR_1[3]),
    .SP(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51779.11-51785.2" *)
  FD1P3IX \storage_1_dat1_reg[3]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(storage_1_TMR_2[3]),
    .Q(storage_1_dat1_TMR_2[3]),
    .SP(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51787.11-51793.2" *)
  FD1P3IX \storage_1_dat1_reg[4]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(storage_1_TMR_0[4]),
    .Q(storage_1_dat1_TMR_0[4]),
    .SP(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51787.11-51793.2" *)
  FD1P3IX \storage_1_dat1_reg[4]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(storage_1_TMR_1[4]),
    .Q(storage_1_dat1_TMR_1[4]),
    .SP(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51787.11-51793.2" *)
  FD1P3IX \storage_1_dat1_reg[4]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(storage_1_TMR_2[4]),
    .Q(storage_1_dat1_TMR_2[4]),
    .SP(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51795.11-51801.2" *)
  FD1P3IX \storage_1_dat1_reg[5]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(storage_1_TMR_0[5]),
    .Q(storage_1_dat1_TMR_0[5]),
    .SP(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51795.11-51801.2" *)
  FD1P3IX \storage_1_dat1_reg[5]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(storage_1_TMR_1[5]),
    .Q(storage_1_dat1_TMR_1[5]),
    .SP(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51795.11-51801.2" *)
  FD1P3IX \storage_1_dat1_reg[5]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(storage_1_TMR_2[5]),
    .Q(storage_1_dat1_TMR_2[5]),
    .SP(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51803.11-51809.2" *)
  FD1P3IX \storage_1_dat1_reg[6]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(storage_1_TMR_0[6]),
    .Q(storage_1_dat1_TMR_0[6]),
    .SP(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51803.11-51809.2" *)
  FD1P3IX \storage_1_dat1_reg[6]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(storage_1_TMR_1[6]),
    .Q(storage_1_dat1_TMR_1[6]),
    .SP(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51803.11-51809.2" *)
  FD1P3IX \storage_1_dat1_reg[6]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(storage_1_TMR_2[6]),
    .Q(storage_1_dat1_TMR_2[6]),
    .SP(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51811.11-51817.2" *)
  FD1P3IX \storage_1_dat1_reg[7]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(storage_1_TMR_0[7]),
    .Q(storage_1_dat1_TMR_0[7]),
    .SP(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51811.11-51817.2" *)
  FD1P3IX \storage_1_dat1_reg[7]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(storage_1_TMR_1[7]),
    .Q(storage_1_dat1_TMR_1[7]),
    .SP(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51811.11-51817.2" *)
  FD1P3IX \storage_1_dat1_reg[7]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(storage_1_TMR_2[7]),
    .Q(storage_1_dat1_TMR_2[7]),
    .SP(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57947.11-57954.2" *)
  DPR16X4 storage_1_ram_0_TMR_0 (
    .DI(main_basesoc_rx_source_payload_data_TMR_0[7:4]),
    .DO(storage_1_TMR_0[7:4]),
    .RAD(main_basesoc_uart_rx_fifo_consume_TMR_0),
    .WAD(main_basesoc_uart_rx_fifo_produce_TMR_0),
    .WCK(sys_clk),
    .WRE(main_basesoc_uart_rx_fifo_wrport_we_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57947.11-57954.2" *)
  DPR16X4 storage_1_ram_0_TMR_1 (
    .DI(main_basesoc_rx_source_payload_data_TMR_1[7:4]),
    .DO(storage_1_TMR_1[7:4]),
    .RAD(main_basesoc_uart_rx_fifo_consume_TMR_1),
    .WAD(main_basesoc_uart_rx_fifo_produce_TMR_1),
    .WCK(sys_clk),
    .WRE(main_basesoc_uart_rx_fifo_wrport_we_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57947.11-57954.2" *)
  DPR16X4 storage_1_ram_0_TMR_2 (
    .DI(main_basesoc_rx_source_payload_data_TMR_2[7:4]),
    .DO(storage_1_TMR_2[7:4]),
    .RAD(main_basesoc_uart_rx_fifo_consume_TMR_2),
    .WAD(main_basesoc_uart_rx_fifo_produce_TMR_2),
    .WCK(sys_clk),
    .WRE(main_basesoc_uart_rx_fifo_wrport_we_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57956.11-57963.2" *)
  DPR16X4 storage_1_ram_TMR_0 (
    .DI(main_basesoc_rx_source_payload_data_TMR_0[3:0]),
    .DO(storage_1_TMR_0[3:0]),
    .RAD(main_basesoc_uart_rx_fifo_consume_TMR_0),
    .WAD(main_basesoc_uart_rx_fifo_produce_TMR_0),
    .WCK(sys_clk),
    .WRE(main_basesoc_uart_rx_fifo_wrport_we_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57956.11-57963.2" *)
  DPR16X4 storage_1_ram_TMR_1 (
    .DI(main_basesoc_rx_source_payload_data_TMR_1[3:0]),
    .DO(storage_1_TMR_1[3:0]),
    .RAD(main_basesoc_uart_rx_fifo_consume_TMR_1),
    .WAD(main_basesoc_uart_rx_fifo_produce_TMR_1),
    .WCK(sys_clk),
    .WRE(main_basesoc_uart_rx_fifo_wrport_we_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57956.11-57963.2" *)
  DPR16X4 storage_1_ram_TMR_2 (
    .DI(main_basesoc_rx_source_payload_data_TMR_2[3:0]),
    .DO(storage_1_TMR_2[3:0]),
    .RAD(main_basesoc_uart_rx_fifo_consume_TMR_2),
    .WAD(main_basesoc_uart_rx_fifo_produce_TMR_2),
    .WCK(sys_clk),
    .WRE(main_basesoc_uart_rx_fifo_wrport_we_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51691.11-51697.2" *)
  FD1P3IX \storage_dat1_reg[0]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(storage_TMR_0[0]),
    .Q(storage_dat1_TMR_0[0]),
    .SP(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51691.11-51697.2" *)
  FD1P3IX \storage_dat1_reg[0]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(storage_TMR_1[0]),
    .Q(storage_dat1_TMR_1[0]),
    .SP(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51691.11-51697.2" *)
  FD1P3IX \storage_dat1_reg[0]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(storage_TMR_2[0]),
    .Q(storage_dat1_TMR_2[0]),
    .SP(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51699.11-51705.2" *)
  FD1P3IX \storage_dat1_reg[1]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(storage_TMR_0[1]),
    .Q(storage_dat1_TMR_0[1]),
    .SP(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51699.11-51705.2" *)
  FD1P3IX \storage_dat1_reg[1]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(storage_TMR_1[1]),
    .Q(storage_dat1_TMR_1[1]),
    .SP(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51699.11-51705.2" *)
  FD1P3IX \storage_dat1_reg[1]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(storage_TMR_2[1]),
    .Q(storage_dat1_TMR_2[1]),
    .SP(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51707.11-51713.2" *)
  FD1P3IX \storage_dat1_reg[2]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(storage_TMR_0[2]),
    .Q(storage_dat1_TMR_0[2]),
    .SP(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51707.11-51713.2" *)
  FD1P3IX \storage_dat1_reg[2]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(storage_TMR_1[2]),
    .Q(storage_dat1_TMR_1[2]),
    .SP(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51707.11-51713.2" *)
  FD1P3IX \storage_dat1_reg[2]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(storage_TMR_2[2]),
    .Q(storage_dat1_TMR_2[2]),
    .SP(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51715.11-51721.2" *)
  FD1P3IX \storage_dat1_reg[3]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(storage_TMR_0[3]),
    .Q(storage_dat1_TMR_0[3]),
    .SP(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51715.11-51721.2" *)
  FD1P3IX \storage_dat1_reg[3]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(storage_TMR_1[3]),
    .Q(storage_dat1_TMR_1[3]),
    .SP(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51715.11-51721.2" *)
  FD1P3IX \storage_dat1_reg[3]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(storage_TMR_2[3]),
    .Q(storage_dat1_TMR_2[3]),
    .SP(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51723.11-51729.2" *)
  FD1P3IX \storage_dat1_reg[4]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(storage_TMR_0[4]),
    .Q(storage_dat1_TMR_0[4]),
    .SP(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51723.11-51729.2" *)
  FD1P3IX \storage_dat1_reg[4]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(storage_TMR_1[4]),
    .Q(storage_dat1_TMR_1[4]),
    .SP(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51723.11-51729.2" *)
  FD1P3IX \storage_dat1_reg[4]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(storage_TMR_2[4]),
    .Q(storage_dat1_TMR_2[4]),
    .SP(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51731.11-51737.2" *)
  FD1P3IX \storage_dat1_reg[5]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(storage_TMR_0[5]),
    .Q(storage_dat1_TMR_0[5]),
    .SP(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51731.11-51737.2" *)
  FD1P3IX \storage_dat1_reg[5]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(storage_TMR_1[5]),
    .Q(storage_dat1_TMR_1[5]),
    .SP(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51731.11-51737.2" *)
  FD1P3IX \storage_dat1_reg[5]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(storage_TMR_2[5]),
    .Q(storage_dat1_TMR_2[5]),
    .SP(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51739.11-51745.2" *)
  FD1P3IX \storage_dat1_reg[6]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(storage_TMR_0[6]),
    .Q(storage_dat1_TMR_0[6]),
    .SP(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51739.11-51745.2" *)
  FD1P3IX \storage_dat1_reg[6]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(storage_TMR_1[6]),
    .Q(storage_dat1_TMR_1[6]),
    .SP(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51739.11-51745.2" *)
  FD1P3IX \storage_dat1_reg[6]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(storage_TMR_2[6]),
    .Q(storage_dat1_TMR_2[6]),
    .SP(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51747.11-51753.2" *)
  FD1P3IX \storage_dat1_reg[7]_TMR_0  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(storage_TMR_0[7]),
    .Q(storage_dat1_TMR_0[7]),
    .SP(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51747.11-51753.2" *)
  FD1P3IX \storage_dat1_reg[7]_TMR_1  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(storage_TMR_1[7]),
    .Q(storage_dat1_TMR_1[7]),
    .SP(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:51747.11-51753.2" *)
  FD1P3IX \storage_dat1_reg[7]_TMR_2  (
    .CD(GND_0),
    .CK(sys_clk),
    .D(storage_TMR_2[7]),
    .Q(storage_dat1_TMR_2[7]),
    .SP(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57965.11-57972.2" *)
  DPR16X4 storage_ram_0_TMR_0 (
    .DI(dsp_join_kb_0_TMR_0[7:4]),
    .DO(storage_TMR_0[7:4]),
    .RAD(main_basesoc_uart_tx_fifo_consume_TMR_0),
    .WAD(main_basesoc_uart_tx_fifo_produce_TMR_0),
    .WCK(sys_clk),
    .WRE(main_basesoc_uart_tx_fifo_wrport_we_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57965.11-57972.2" *)
  DPR16X4 storage_ram_0_TMR_1 (
    .DI(dsp_join_kb_0_TMR_1[7:4]),
    .DO(storage_TMR_1[7:4]),
    .RAD(main_basesoc_uart_tx_fifo_consume_TMR_1),
    .WAD(main_basesoc_uart_tx_fifo_produce_TMR_1),
    .WCK(sys_clk),
    .WRE(main_basesoc_uart_tx_fifo_wrport_we_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57965.11-57972.2" *)
  DPR16X4 storage_ram_0_TMR_2 (
    .DI(dsp_join_kb_0_TMR_2[7:4]),
    .DO(storage_TMR_2[7:4]),
    .RAD(main_basesoc_uart_tx_fifo_consume_TMR_2),
    .WAD(main_basesoc_uart_tx_fifo_produce_TMR_2),
    .WCK(sys_clk),
    .WRE(main_basesoc_uart_tx_fifo_wrport_we_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57974.11-57981.2" *)
  DPR16X4 storage_ram_TMR_0 (
    .DI(dsp_join_kb_0_TMR_0[3:0]),
    .DO(storage_TMR_0[3:0]),
    .RAD(main_basesoc_uart_tx_fifo_consume_TMR_0),
    .WAD(main_basesoc_uart_tx_fifo_produce_TMR_0),
    .WCK(sys_clk),
    .WRE(main_basesoc_uart_tx_fifo_wrport_we_TMR_0)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57974.11-57981.2" *)
  DPR16X4 storage_ram_TMR_1 (
    .DI(dsp_join_kb_0_TMR_1[3:0]),
    .DO(storage_TMR_1[3:0]),
    .RAD(main_basesoc_uart_tx_fifo_consume_TMR_1),
    .WAD(main_basesoc_uart_tx_fifo_produce_TMR_1),
    .WCK(sys_clk),
    .WRE(main_basesoc_uart_tx_fifo_wrport_we_TMR_1)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57974.11-57981.2" *)
  DPR16X4 storage_ram_TMR_2 (
    .DI(dsp_join_kb_0_TMR_2[3:0]),
    .DO(storage_TMR_2[3:0]),
    .RAD(main_basesoc_uart_tx_fifo_consume_TMR_2),
    .WAD(main_basesoc_uart_tx_fifo_produce_TMR_2),
    .WCK(sys_clk),
    .WRE(main_basesoc_uart_tx_fifo_wrport_we_TMR_2)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56746.8-56759.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_cry_0_0_TMR_0 (
    .A0(VCC_TMR_0),
    .A1(un1_main_basesoc_bus_errors_1_0_TMR_0[0]),
    .B0(main_basesoc_bus_errors_0_sqmuxa_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(GND_0),
    .COUT(un1_main_basesoc_bus_errors_1_cry_0_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un1_main_basesoc_bus_errors_1_cry_0_0_S0_TMR_0),
    .S1(un1_main_basesoc_bus_errors_1_TMR_0[0])
  );
  defparam un1_main_basesoc_bus_errors_1_cry_0_0_TMR_0.INIT0 = "50CC";
  defparam un1_main_basesoc_bus_errors_1_cry_0_0_TMR_0.INIT1 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_0_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56746.8-56759.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_cry_0_0_TMR_1 (
    .A0(VCC_TMR_1),
    .A1(un1_main_basesoc_bus_errors_1_0_TMR_1[0]),
    .B0(main_basesoc_bus_errors_0_sqmuxa_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(GND_0),
    .COUT(un1_main_basesoc_bus_errors_1_cry_0_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un1_main_basesoc_bus_errors_1_cry_0_0_S0_TMR_1),
    .S1(un1_main_basesoc_bus_errors_1_TMR_1[0])
  );
  defparam un1_main_basesoc_bus_errors_1_cry_0_0_TMR_1.INIT0 = "50CC";
  defparam un1_main_basesoc_bus_errors_1_cry_0_0_TMR_1.INIT1 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_0_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56746.8-56759.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_cry_0_0_TMR_2 (
    .A0(VCC_TMR_2),
    .A1(un1_main_basesoc_bus_errors_1_0_TMR_2[0]),
    .B0(main_basesoc_bus_errors_0_sqmuxa_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(GND_0),
    .COUT(un1_main_basesoc_bus_errors_1_cry_0_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un1_main_basesoc_bus_errors_1_cry_0_0_S0_TMR_2),
    .S1(un1_main_basesoc_bus_errors_1_TMR_2[0])
  );
  defparam un1_main_basesoc_bus_errors_1_cry_0_0_TMR_2.INIT0 = "50CC";
  defparam un1_main_basesoc_bus_errors_1_cry_0_0_TMR_2.INIT1 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_0_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56639.8-56652.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_cry_11_0_TMR_0 (
    .A0(un1_main_basesoc_bus_errors_1_0_TMR_0[11]),
    .A1(un1_main_basesoc_bus_errors_1_0_TMR_0[12]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(un1_main_basesoc_bus_errors_1_cry_10_TMR_0),
    .COUT(un1_main_basesoc_bus_errors_1_cry_12_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un1_main_basesoc_bus_errors_1_TMR_0[11]),
    .S1(un1_main_basesoc_bus_errors_1_TMR_0[12])
  );
  defparam un1_main_basesoc_bus_errors_1_cry_11_0_TMR_0.INIT0 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_11_0_TMR_0.INIT1 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_11_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56639.8-56652.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_cry_11_0_TMR_1 (
    .A0(un1_main_basesoc_bus_errors_1_0_TMR_1[11]),
    .A1(un1_main_basesoc_bus_errors_1_0_TMR_1[12]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(un1_main_basesoc_bus_errors_1_cry_10_TMR_1),
    .COUT(un1_main_basesoc_bus_errors_1_cry_12_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un1_main_basesoc_bus_errors_1_TMR_1[11]),
    .S1(un1_main_basesoc_bus_errors_1_TMR_1[12])
  );
  defparam un1_main_basesoc_bus_errors_1_cry_11_0_TMR_1.INIT0 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_11_0_TMR_1.INIT1 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_11_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56639.8-56652.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_cry_11_0_TMR_2 (
    .A0(un1_main_basesoc_bus_errors_1_0_TMR_2[11]),
    .A1(un1_main_basesoc_bus_errors_1_0_TMR_2[12]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(un1_main_basesoc_bus_errors_1_cry_10_TMR_2),
    .COUT(un1_main_basesoc_bus_errors_1_cry_12_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un1_main_basesoc_bus_errors_1_TMR_2[11]),
    .S1(un1_main_basesoc_bus_errors_1_TMR_2[12])
  );
  defparam un1_main_basesoc_bus_errors_1_cry_11_0_TMR_2.INIT0 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_11_0_TMR_2.INIT1 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_11_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56621.8-56634.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_cry_13_0_TMR_0 (
    .A0(un1_main_basesoc_bus_errors_1_0_TMR_0[13]),
    .A1(un1_main_basesoc_bus_errors_1_0_TMR_0[14]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(un1_main_basesoc_bus_errors_1_cry_12_TMR_0),
    .COUT(un1_main_basesoc_bus_errors_1_cry_14_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un1_main_basesoc_bus_errors_1_TMR_0[13]),
    .S1(un1_main_basesoc_bus_errors_1_TMR_0[14])
  );
  defparam un1_main_basesoc_bus_errors_1_cry_13_0_TMR_0.INIT0 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_13_0_TMR_0.INIT1 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_13_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56621.8-56634.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_cry_13_0_TMR_1 (
    .A0(un1_main_basesoc_bus_errors_1_0_TMR_1[13]),
    .A1(un1_main_basesoc_bus_errors_1_0_TMR_1[14]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(un1_main_basesoc_bus_errors_1_cry_12_TMR_1),
    .COUT(un1_main_basesoc_bus_errors_1_cry_14_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un1_main_basesoc_bus_errors_1_TMR_1[13]),
    .S1(un1_main_basesoc_bus_errors_1_TMR_1[14])
  );
  defparam un1_main_basesoc_bus_errors_1_cry_13_0_TMR_1.INIT0 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_13_0_TMR_1.INIT1 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_13_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56621.8-56634.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_cry_13_0_TMR_2 (
    .A0(un1_main_basesoc_bus_errors_1_0_TMR_2[13]),
    .A1(un1_main_basesoc_bus_errors_1_0_TMR_2[14]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(un1_main_basesoc_bus_errors_1_cry_12_TMR_2),
    .COUT(un1_main_basesoc_bus_errors_1_cry_14_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un1_main_basesoc_bus_errors_1_TMR_2[13]),
    .S1(un1_main_basesoc_bus_errors_1_TMR_2[14])
  );
  defparam un1_main_basesoc_bus_errors_1_cry_13_0_TMR_2.INIT0 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_13_0_TMR_2.INIT1 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_13_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56603.8-56616.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_cry_15_0_TMR_0 (
    .A0(un1_main_basesoc_bus_errors_1_0_TMR_0[15]),
    .A1(un1_main_basesoc_bus_errors_1_0_TMR_0[16]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(un1_main_basesoc_bus_errors_1_cry_14_TMR_0),
    .COUT(un1_main_basesoc_bus_errors_1_cry_16_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un1_main_basesoc_bus_errors_1_TMR_0[15]),
    .S1(un1_main_basesoc_bus_errors_1_TMR_0[16])
  );
  defparam un1_main_basesoc_bus_errors_1_cry_15_0_TMR_0.INIT0 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_15_0_TMR_0.INIT1 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_15_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56603.8-56616.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_cry_15_0_TMR_1 (
    .A0(un1_main_basesoc_bus_errors_1_0_TMR_1[15]),
    .A1(un1_main_basesoc_bus_errors_1_0_TMR_1[16]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(un1_main_basesoc_bus_errors_1_cry_14_TMR_1),
    .COUT(un1_main_basesoc_bus_errors_1_cry_16_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un1_main_basesoc_bus_errors_1_TMR_1[15]),
    .S1(un1_main_basesoc_bus_errors_1_TMR_1[16])
  );
  defparam un1_main_basesoc_bus_errors_1_cry_15_0_TMR_1.INIT0 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_15_0_TMR_1.INIT1 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_15_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56603.8-56616.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_cry_15_0_TMR_2 (
    .A0(un1_main_basesoc_bus_errors_1_0_TMR_2[15]),
    .A1(un1_main_basesoc_bus_errors_1_0_TMR_2[16]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(un1_main_basesoc_bus_errors_1_cry_14_TMR_2),
    .COUT(un1_main_basesoc_bus_errors_1_cry_16_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un1_main_basesoc_bus_errors_1_TMR_2[15]),
    .S1(un1_main_basesoc_bus_errors_1_TMR_2[16])
  );
  defparam un1_main_basesoc_bus_errors_1_cry_15_0_TMR_2.INIT0 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_15_0_TMR_2.INIT1 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_15_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56585.8-56598.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_cry_17_0_TMR_0 (
    .A0(un1_main_basesoc_bus_errors_1_0_TMR_0[17]),
    .A1(un1_main_basesoc_bus_errors_1_0_TMR_0[18]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(un1_main_basesoc_bus_errors_1_cry_16_TMR_0),
    .COUT(un1_main_basesoc_bus_errors_1_cry_18_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un1_main_basesoc_bus_errors_1_TMR_0[17]),
    .S1(un1_main_basesoc_bus_errors_1_TMR_0[18])
  );
  defparam un1_main_basesoc_bus_errors_1_cry_17_0_TMR_0.INIT0 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_17_0_TMR_0.INIT1 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_17_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56585.8-56598.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_cry_17_0_TMR_1 (
    .A0(un1_main_basesoc_bus_errors_1_0_TMR_1[17]),
    .A1(un1_main_basesoc_bus_errors_1_0_TMR_1[18]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(un1_main_basesoc_bus_errors_1_cry_16_TMR_1),
    .COUT(un1_main_basesoc_bus_errors_1_cry_18_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un1_main_basesoc_bus_errors_1_TMR_1[17]),
    .S1(un1_main_basesoc_bus_errors_1_TMR_1[18])
  );
  defparam un1_main_basesoc_bus_errors_1_cry_17_0_TMR_1.INIT0 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_17_0_TMR_1.INIT1 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_17_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56585.8-56598.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_cry_17_0_TMR_2 (
    .A0(un1_main_basesoc_bus_errors_1_0_TMR_2[17]),
    .A1(un1_main_basesoc_bus_errors_1_0_TMR_2[18]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(un1_main_basesoc_bus_errors_1_cry_16_TMR_2),
    .COUT(un1_main_basesoc_bus_errors_1_cry_18_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un1_main_basesoc_bus_errors_1_TMR_2[17]),
    .S1(un1_main_basesoc_bus_errors_1_TMR_2[18])
  );
  defparam un1_main_basesoc_bus_errors_1_cry_17_0_TMR_2.INIT0 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_17_0_TMR_2.INIT1 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_17_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56567.8-56580.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_cry_19_0_TMR_0 (
    .A0(un1_main_basesoc_bus_errors_1_0_TMR_0[19]),
    .A1(un1_main_basesoc_bus_errors_1_0_TMR_0[20]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(un1_main_basesoc_bus_errors_1_cry_18_TMR_0),
    .COUT(un1_main_basesoc_bus_errors_1_cry_20_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un1_main_basesoc_bus_errors_1_TMR_0[19]),
    .S1(un1_main_basesoc_bus_errors_1_TMR_0[20])
  );
  defparam un1_main_basesoc_bus_errors_1_cry_19_0_TMR_0.INIT0 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_19_0_TMR_0.INIT1 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_19_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56567.8-56580.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_cry_19_0_TMR_1 (
    .A0(un1_main_basesoc_bus_errors_1_0_TMR_1[19]),
    .A1(un1_main_basesoc_bus_errors_1_0_TMR_1[20]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(un1_main_basesoc_bus_errors_1_cry_18_TMR_1),
    .COUT(un1_main_basesoc_bus_errors_1_cry_20_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un1_main_basesoc_bus_errors_1_TMR_1[19]),
    .S1(un1_main_basesoc_bus_errors_1_TMR_1[20])
  );
  defparam un1_main_basesoc_bus_errors_1_cry_19_0_TMR_1.INIT0 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_19_0_TMR_1.INIT1 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_19_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56567.8-56580.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_cry_19_0_TMR_2 (
    .A0(un1_main_basesoc_bus_errors_1_0_TMR_2[19]),
    .A1(un1_main_basesoc_bus_errors_1_0_TMR_2[20]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(un1_main_basesoc_bus_errors_1_cry_18_TMR_2),
    .COUT(un1_main_basesoc_bus_errors_1_cry_20_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un1_main_basesoc_bus_errors_1_TMR_2[19]),
    .S1(un1_main_basesoc_bus_errors_1_TMR_2[20])
  );
  defparam un1_main_basesoc_bus_errors_1_cry_19_0_TMR_2.INIT0 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_19_0_TMR_2.INIT1 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_19_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56729.8-56742.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_cry_1_0_TMR_0 (
    .A0(un1_main_basesoc_bus_errors_1_0_TMR_0[1]),
    .A1(un1_main_basesoc_bus_errors_1_0_TMR_0[2]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(un1_main_basesoc_bus_errors_1_cry_0_TMR_0),
    .COUT(un1_main_basesoc_bus_errors_1_cry_2_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un1_main_basesoc_bus_errors_1_TMR_0[1]),
    .S1(un1_main_basesoc_bus_errors_1_TMR_0[2])
  );
  defparam un1_main_basesoc_bus_errors_1_cry_1_0_TMR_0.INIT0 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_1_0_TMR_0.INIT1 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_1_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56729.8-56742.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_cry_1_0_TMR_1 (
    .A0(un1_main_basesoc_bus_errors_1_0_TMR_1[1]),
    .A1(un1_main_basesoc_bus_errors_1_0_TMR_1[2]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(un1_main_basesoc_bus_errors_1_cry_0_TMR_1),
    .COUT(un1_main_basesoc_bus_errors_1_cry_2_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un1_main_basesoc_bus_errors_1_TMR_1[1]),
    .S1(un1_main_basesoc_bus_errors_1_TMR_1[2])
  );
  defparam un1_main_basesoc_bus_errors_1_cry_1_0_TMR_1.INIT0 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_1_0_TMR_1.INIT1 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_1_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56729.8-56742.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_cry_1_0_TMR_2 (
    .A0(un1_main_basesoc_bus_errors_1_0_TMR_2[1]),
    .A1(un1_main_basesoc_bus_errors_1_0_TMR_2[2]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(un1_main_basesoc_bus_errors_1_cry_0_TMR_2),
    .COUT(un1_main_basesoc_bus_errors_1_cry_2_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un1_main_basesoc_bus_errors_1_TMR_2[1]),
    .S1(un1_main_basesoc_bus_errors_1_TMR_2[2])
  );
  defparam un1_main_basesoc_bus_errors_1_cry_1_0_TMR_2.INIT0 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_1_0_TMR_2.INIT1 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_1_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56549.8-56562.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_cry_21_0_TMR_0 (
    .A0(un1_main_basesoc_bus_errors_1_0_TMR_0[21]),
    .A1(un1_main_basesoc_bus_errors_1_0_TMR_0[22]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(un1_main_basesoc_bus_errors_1_cry_20_TMR_0),
    .COUT(un1_main_basesoc_bus_errors_1_cry_22_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un1_main_basesoc_bus_errors_1_TMR_0[21]),
    .S1(un1_main_basesoc_bus_errors_1_TMR_0[22])
  );
  defparam un1_main_basesoc_bus_errors_1_cry_21_0_TMR_0.INIT0 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_21_0_TMR_0.INIT1 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_21_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56549.8-56562.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_cry_21_0_TMR_1 (
    .A0(un1_main_basesoc_bus_errors_1_0_TMR_1[21]),
    .A1(un1_main_basesoc_bus_errors_1_0_TMR_1[22]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(un1_main_basesoc_bus_errors_1_cry_20_TMR_1),
    .COUT(un1_main_basesoc_bus_errors_1_cry_22_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un1_main_basesoc_bus_errors_1_TMR_1[21]),
    .S1(un1_main_basesoc_bus_errors_1_TMR_1[22])
  );
  defparam un1_main_basesoc_bus_errors_1_cry_21_0_TMR_1.INIT0 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_21_0_TMR_1.INIT1 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_21_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56549.8-56562.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_cry_21_0_TMR_2 (
    .A0(un1_main_basesoc_bus_errors_1_0_TMR_2[21]),
    .A1(un1_main_basesoc_bus_errors_1_0_TMR_2[22]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(un1_main_basesoc_bus_errors_1_cry_20_TMR_2),
    .COUT(un1_main_basesoc_bus_errors_1_cry_22_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un1_main_basesoc_bus_errors_1_TMR_2[21]),
    .S1(un1_main_basesoc_bus_errors_1_TMR_2[22])
  );
  defparam un1_main_basesoc_bus_errors_1_cry_21_0_TMR_2.INIT0 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_21_0_TMR_2.INIT1 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_21_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56531.8-56544.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_cry_23_0_TMR_0 (
    .A0(un1_main_basesoc_bus_errors_1_0_TMR_0[23]),
    .A1(un1_main_basesoc_bus_errors_1_0_TMR_0[24]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(un1_main_basesoc_bus_errors_1_cry_22_TMR_0),
    .COUT(un1_main_basesoc_bus_errors_1_cry_24_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un1_main_basesoc_bus_errors_1_TMR_0[23]),
    .S1(un1_main_basesoc_bus_errors_1_TMR_0[24])
  );
  defparam un1_main_basesoc_bus_errors_1_cry_23_0_TMR_0.INIT0 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_23_0_TMR_0.INIT1 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_23_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56531.8-56544.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_cry_23_0_TMR_1 (
    .A0(un1_main_basesoc_bus_errors_1_0_TMR_1[23]),
    .A1(un1_main_basesoc_bus_errors_1_0_TMR_1[24]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(un1_main_basesoc_bus_errors_1_cry_22_TMR_1),
    .COUT(un1_main_basesoc_bus_errors_1_cry_24_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un1_main_basesoc_bus_errors_1_TMR_1[23]),
    .S1(un1_main_basesoc_bus_errors_1_TMR_1[24])
  );
  defparam un1_main_basesoc_bus_errors_1_cry_23_0_TMR_1.INIT0 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_23_0_TMR_1.INIT1 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_23_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56531.8-56544.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_cry_23_0_TMR_2 (
    .A0(un1_main_basesoc_bus_errors_1_0_TMR_2[23]),
    .A1(un1_main_basesoc_bus_errors_1_0_TMR_2[24]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(un1_main_basesoc_bus_errors_1_cry_22_TMR_2),
    .COUT(un1_main_basesoc_bus_errors_1_cry_24_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un1_main_basesoc_bus_errors_1_TMR_2[23]),
    .S1(un1_main_basesoc_bus_errors_1_TMR_2[24])
  );
  defparam un1_main_basesoc_bus_errors_1_cry_23_0_TMR_2.INIT0 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_23_0_TMR_2.INIT1 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_23_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56513.8-56526.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_cry_25_0_TMR_0 (
    .A0(un1_main_basesoc_bus_errors_1_0_TMR_0[25]),
    .A1(un1_main_basesoc_bus_errors_1_0_TMR_0[26]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(un1_main_basesoc_bus_errors_1_cry_24_TMR_0),
    .COUT(un1_main_basesoc_bus_errors_1_cry_26_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un1_main_basesoc_bus_errors_1_TMR_0[25]),
    .S1(un1_main_basesoc_bus_errors_1_TMR_0[26])
  );
  defparam un1_main_basesoc_bus_errors_1_cry_25_0_TMR_0.INIT0 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_25_0_TMR_0.INIT1 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_25_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56513.8-56526.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_cry_25_0_TMR_1 (
    .A0(un1_main_basesoc_bus_errors_1_0_TMR_1[25]),
    .A1(un1_main_basesoc_bus_errors_1_0_TMR_1[26]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(un1_main_basesoc_bus_errors_1_cry_24_TMR_1),
    .COUT(un1_main_basesoc_bus_errors_1_cry_26_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un1_main_basesoc_bus_errors_1_TMR_1[25]),
    .S1(un1_main_basesoc_bus_errors_1_TMR_1[26])
  );
  defparam un1_main_basesoc_bus_errors_1_cry_25_0_TMR_1.INIT0 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_25_0_TMR_1.INIT1 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_25_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56513.8-56526.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_cry_25_0_TMR_2 (
    .A0(un1_main_basesoc_bus_errors_1_0_TMR_2[25]),
    .A1(un1_main_basesoc_bus_errors_1_0_TMR_2[26]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(un1_main_basesoc_bus_errors_1_cry_24_TMR_2),
    .COUT(un1_main_basesoc_bus_errors_1_cry_26_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un1_main_basesoc_bus_errors_1_TMR_2[25]),
    .S1(un1_main_basesoc_bus_errors_1_TMR_2[26])
  );
  defparam un1_main_basesoc_bus_errors_1_cry_25_0_TMR_2.INIT0 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_25_0_TMR_2.INIT1 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_25_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56495.8-56508.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_cry_27_0_TMR_0 (
    .A0(un1_main_basesoc_bus_errors_1_0_TMR_0[27]),
    .A1(un1_main_basesoc_bus_errors_1_0_TMR_0[28]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(un1_main_basesoc_bus_errors_1_cry_26_TMR_0),
    .COUT(un1_main_basesoc_bus_errors_1_cry_28_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un1_main_basesoc_bus_errors_1_TMR_0[27]),
    .S1(un1_main_basesoc_bus_errors_1_TMR_0[28])
  );
  defparam un1_main_basesoc_bus_errors_1_cry_27_0_TMR_0.INIT0 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_27_0_TMR_0.INIT1 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_27_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56495.8-56508.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_cry_27_0_TMR_1 (
    .A0(un1_main_basesoc_bus_errors_1_0_TMR_1[27]),
    .A1(un1_main_basesoc_bus_errors_1_0_TMR_1[28]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(un1_main_basesoc_bus_errors_1_cry_26_TMR_1),
    .COUT(un1_main_basesoc_bus_errors_1_cry_28_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un1_main_basesoc_bus_errors_1_TMR_1[27]),
    .S1(un1_main_basesoc_bus_errors_1_TMR_1[28])
  );
  defparam un1_main_basesoc_bus_errors_1_cry_27_0_TMR_1.INIT0 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_27_0_TMR_1.INIT1 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_27_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56495.8-56508.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_cry_27_0_TMR_2 (
    .A0(un1_main_basesoc_bus_errors_1_0_TMR_2[27]),
    .A1(un1_main_basesoc_bus_errors_1_0_TMR_2[28]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(un1_main_basesoc_bus_errors_1_cry_26_TMR_2),
    .COUT(un1_main_basesoc_bus_errors_1_cry_28_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un1_main_basesoc_bus_errors_1_TMR_2[27]),
    .S1(un1_main_basesoc_bus_errors_1_TMR_2[28])
  );
  defparam un1_main_basesoc_bus_errors_1_cry_27_0_TMR_2.INIT0 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_27_0_TMR_2.INIT1 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_27_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56477.8-56490.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_cry_29_0_TMR_0 (
    .A0(un1_main_basesoc_bus_errors_1_0_TMR_0[29]),
    .A1(un1_main_basesoc_bus_errors_1_0_TMR_0[30]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(un1_main_basesoc_bus_errors_1_cry_28_TMR_0),
    .COUT(un1_main_basesoc_bus_errors_1_cry_30_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un1_main_basesoc_bus_errors_1_TMR_0[29]),
    .S1(un1_main_basesoc_bus_errors_1_TMR_0[30])
  );
  defparam un1_main_basesoc_bus_errors_1_cry_29_0_TMR_0.INIT0 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_29_0_TMR_0.INIT1 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_29_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56477.8-56490.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_cry_29_0_TMR_1 (
    .A0(un1_main_basesoc_bus_errors_1_0_TMR_1[29]),
    .A1(un1_main_basesoc_bus_errors_1_0_TMR_1[30]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(un1_main_basesoc_bus_errors_1_cry_28_TMR_1),
    .COUT(un1_main_basesoc_bus_errors_1_cry_30_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un1_main_basesoc_bus_errors_1_TMR_1[29]),
    .S1(un1_main_basesoc_bus_errors_1_TMR_1[30])
  );
  defparam un1_main_basesoc_bus_errors_1_cry_29_0_TMR_1.INIT0 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_29_0_TMR_1.INIT1 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_29_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56477.8-56490.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_cry_29_0_TMR_2 (
    .A0(un1_main_basesoc_bus_errors_1_0_TMR_2[29]),
    .A1(un1_main_basesoc_bus_errors_1_0_TMR_2[30]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(un1_main_basesoc_bus_errors_1_cry_28_TMR_2),
    .COUT(un1_main_basesoc_bus_errors_1_cry_30_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un1_main_basesoc_bus_errors_1_TMR_2[29]),
    .S1(un1_main_basesoc_bus_errors_1_TMR_2[30])
  );
  defparam un1_main_basesoc_bus_errors_1_cry_29_0_TMR_2.INIT0 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_29_0_TMR_2.INIT1 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_29_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56711.8-56724.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_cry_3_0_TMR_0 (
    .A0(un1_main_basesoc_bus_errors_1_0_TMR_0[3]),
    .A1(un1_main_basesoc_bus_errors_1_0_TMR_0[4]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(un1_main_basesoc_bus_errors_1_cry_2_TMR_0),
    .COUT(un1_main_basesoc_bus_errors_1_cry_4_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un1_main_basesoc_bus_errors_1_TMR_0[3]),
    .S1(un1_main_basesoc_bus_errors_1_TMR_0[4])
  );
  defparam un1_main_basesoc_bus_errors_1_cry_3_0_TMR_0.INIT0 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_3_0_TMR_0.INIT1 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_3_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56711.8-56724.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_cry_3_0_TMR_1 (
    .A0(un1_main_basesoc_bus_errors_1_0_TMR_1[3]),
    .A1(un1_main_basesoc_bus_errors_1_0_TMR_1[4]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(un1_main_basesoc_bus_errors_1_cry_2_TMR_1),
    .COUT(un1_main_basesoc_bus_errors_1_cry_4_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un1_main_basesoc_bus_errors_1_TMR_1[3]),
    .S1(un1_main_basesoc_bus_errors_1_TMR_1[4])
  );
  defparam un1_main_basesoc_bus_errors_1_cry_3_0_TMR_1.INIT0 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_3_0_TMR_1.INIT1 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_3_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56711.8-56724.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_cry_3_0_TMR_2 (
    .A0(un1_main_basesoc_bus_errors_1_0_TMR_2[3]),
    .A1(un1_main_basesoc_bus_errors_1_0_TMR_2[4]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(un1_main_basesoc_bus_errors_1_cry_2_TMR_2),
    .COUT(un1_main_basesoc_bus_errors_1_cry_4_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un1_main_basesoc_bus_errors_1_TMR_2[3]),
    .S1(un1_main_basesoc_bus_errors_1_TMR_2[4])
  );
  defparam un1_main_basesoc_bus_errors_1_cry_3_0_TMR_2.INIT0 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_3_0_TMR_2.INIT1 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_3_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56693.8-56706.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_cry_5_0_TMR_0 (
    .A0(un1_main_basesoc_bus_errors_1_0_TMR_0[5]),
    .A1(un1_main_basesoc_bus_errors_1_0_TMR_0[6]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(un1_main_basesoc_bus_errors_1_cry_4_TMR_0),
    .COUT(un1_main_basesoc_bus_errors_1_cry_6_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un1_main_basesoc_bus_errors_1_TMR_0[5]),
    .S1(un1_main_basesoc_bus_errors_1_TMR_0[6])
  );
  defparam un1_main_basesoc_bus_errors_1_cry_5_0_TMR_0.INIT0 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_5_0_TMR_0.INIT1 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_5_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56693.8-56706.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_cry_5_0_TMR_1 (
    .A0(un1_main_basesoc_bus_errors_1_0_TMR_1[5]),
    .A1(un1_main_basesoc_bus_errors_1_0_TMR_1[6]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(un1_main_basesoc_bus_errors_1_cry_4_TMR_1),
    .COUT(un1_main_basesoc_bus_errors_1_cry_6_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un1_main_basesoc_bus_errors_1_TMR_1[5]),
    .S1(un1_main_basesoc_bus_errors_1_TMR_1[6])
  );
  defparam un1_main_basesoc_bus_errors_1_cry_5_0_TMR_1.INIT0 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_5_0_TMR_1.INIT1 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_5_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56693.8-56706.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_cry_5_0_TMR_2 (
    .A0(un1_main_basesoc_bus_errors_1_0_TMR_2[5]),
    .A1(un1_main_basesoc_bus_errors_1_0_TMR_2[6]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(un1_main_basesoc_bus_errors_1_cry_4_TMR_2),
    .COUT(un1_main_basesoc_bus_errors_1_cry_6_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un1_main_basesoc_bus_errors_1_TMR_2[5]),
    .S1(un1_main_basesoc_bus_errors_1_TMR_2[6])
  );
  defparam un1_main_basesoc_bus_errors_1_cry_5_0_TMR_2.INIT0 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_5_0_TMR_2.INIT1 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_5_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56675.8-56688.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_cry_7_0_TMR_0 (
    .A0(un1_main_basesoc_bus_errors_1_0_TMR_0[7]),
    .A1(un1_main_basesoc_bus_errors_1_0_TMR_0[8]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(un1_main_basesoc_bus_errors_1_cry_6_TMR_0),
    .COUT(un1_main_basesoc_bus_errors_1_cry_8_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un1_main_basesoc_bus_errors_1_TMR_0[7]),
    .S1(un1_main_basesoc_bus_errors_1_TMR_0[8])
  );
  defparam un1_main_basesoc_bus_errors_1_cry_7_0_TMR_0.INIT0 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_7_0_TMR_0.INIT1 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_7_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56675.8-56688.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_cry_7_0_TMR_1 (
    .A0(un1_main_basesoc_bus_errors_1_0_TMR_1[7]),
    .A1(un1_main_basesoc_bus_errors_1_0_TMR_1[8]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(un1_main_basesoc_bus_errors_1_cry_6_TMR_1),
    .COUT(un1_main_basesoc_bus_errors_1_cry_8_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un1_main_basesoc_bus_errors_1_TMR_1[7]),
    .S1(un1_main_basesoc_bus_errors_1_TMR_1[8])
  );
  defparam un1_main_basesoc_bus_errors_1_cry_7_0_TMR_1.INIT0 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_7_0_TMR_1.INIT1 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_7_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56675.8-56688.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_cry_7_0_TMR_2 (
    .A0(un1_main_basesoc_bus_errors_1_0_TMR_2[7]),
    .A1(un1_main_basesoc_bus_errors_1_0_TMR_2[8]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(un1_main_basesoc_bus_errors_1_cry_6_TMR_2),
    .COUT(un1_main_basesoc_bus_errors_1_cry_8_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un1_main_basesoc_bus_errors_1_TMR_2[7]),
    .S1(un1_main_basesoc_bus_errors_1_TMR_2[8])
  );
  defparam un1_main_basesoc_bus_errors_1_cry_7_0_TMR_2.INIT0 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_7_0_TMR_2.INIT1 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_7_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56657.8-56670.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_cry_9_0_TMR_0 (
    .A0(un1_main_basesoc_bus_errors_1_0_TMR_0[9]),
    .A1(un1_main_basesoc_bus_errors_1_0_TMR_0[10]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(un1_main_basesoc_bus_errors_1_cry_8_TMR_0),
    .COUT(un1_main_basesoc_bus_errors_1_cry_10_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un1_main_basesoc_bus_errors_1_TMR_0[9]),
    .S1(un1_main_basesoc_bus_errors_1_TMR_0[10])
  );
  defparam un1_main_basesoc_bus_errors_1_cry_9_0_TMR_0.INIT0 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_9_0_TMR_0.INIT1 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_9_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56657.8-56670.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_cry_9_0_TMR_1 (
    .A0(un1_main_basesoc_bus_errors_1_0_TMR_1[9]),
    .A1(un1_main_basesoc_bus_errors_1_0_TMR_1[10]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(un1_main_basesoc_bus_errors_1_cry_8_TMR_1),
    .COUT(un1_main_basesoc_bus_errors_1_cry_10_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un1_main_basesoc_bus_errors_1_TMR_1[9]),
    .S1(un1_main_basesoc_bus_errors_1_TMR_1[10])
  );
  defparam un1_main_basesoc_bus_errors_1_cry_9_0_TMR_1.INIT0 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_9_0_TMR_1.INIT1 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_9_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56657.8-56670.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_cry_9_0_TMR_2 (
    .A0(un1_main_basesoc_bus_errors_1_0_TMR_2[9]),
    .A1(un1_main_basesoc_bus_errors_1_0_TMR_2[10]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(un1_main_basesoc_bus_errors_1_cry_8_TMR_2),
    .COUT(un1_main_basesoc_bus_errors_1_cry_10_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un1_main_basesoc_bus_errors_1_TMR_2[9]),
    .S1(un1_main_basesoc_bus_errors_1_TMR_2[10])
  );
  defparam un1_main_basesoc_bus_errors_1_cry_9_0_TMR_2.INIT0 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_9_0_TMR_2.INIT1 = "A033";
  defparam un1_main_basesoc_bus_errors_1_cry_9_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56459.8-56472.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_s_31_0_TMR_0 (
    .A0(un1_main_basesoc_bus_errors_1_0_TMR_0[31]),
    .A1(VCC_TMR_0),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(un1_main_basesoc_bus_errors_1_cry_30_TMR_0),
    .COUT(un1_main_basesoc_bus_errors_1_s_31_0_COUT_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un1_main_basesoc_bus_errors_1_TMR_0[31]),
    .S1(un1_main_basesoc_bus_errors_1_s_31_0_S1_TMR_0)
  );
  defparam un1_main_basesoc_bus_errors_1_s_31_0_TMR_0.INIT0 = "A033";
  defparam un1_main_basesoc_bus_errors_1_s_31_0_TMR_0.INIT1 = "5033";
  defparam un1_main_basesoc_bus_errors_1_s_31_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56459.8-56472.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_s_31_0_TMR_1 (
    .A0(un1_main_basesoc_bus_errors_1_0_TMR_1[31]),
    .A1(VCC_TMR_1),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(un1_main_basesoc_bus_errors_1_cry_30_TMR_1),
    .COUT(un1_main_basesoc_bus_errors_1_s_31_0_COUT_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un1_main_basesoc_bus_errors_1_TMR_1[31]),
    .S1(un1_main_basesoc_bus_errors_1_s_31_0_S1_TMR_1)
  );
  defparam un1_main_basesoc_bus_errors_1_s_31_0_TMR_1.INIT0 = "A033";
  defparam un1_main_basesoc_bus_errors_1_s_31_0_TMR_1.INIT1 = "5033";
  defparam un1_main_basesoc_bus_errors_1_s_31_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56459.8-56472.2" *)
  CCU2 un1_main_basesoc_bus_errors_1_s_31_0_TMR_2 (
    .A0(un1_main_basesoc_bus_errors_1_0_TMR_2[31]),
    .A1(VCC_TMR_2),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(un1_main_basesoc_bus_errors_1_cry_30_TMR_2),
    .COUT(un1_main_basesoc_bus_errors_1_s_31_0_COUT_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un1_main_basesoc_bus_errors_1_TMR_2[31]),
    .S1(un1_main_basesoc_bus_errors_1_s_31_0_S1_TMR_2)
  );
  defparam un1_main_basesoc_bus_errors_1_s_31_0_TMR_2.INIT0 = "A033";
  defparam un1_main_basesoc_bus_errors_1_s_31_0_TMR_2.INIT1 = "5033";
  defparam un1_main_basesoc_bus_errors_1_s_31_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55826.8-55832.2" *)
  LUT4 un1_main_basesoc_uart_rx_fifo_consume_ac0_1_TMR_0 (
    .A(main_basesoc_uart_rx_fifo_consume_TMR_0[0]),
    .B(main_basesoc_uart_rx_fifo_consume_TMR_0[1]),
    .C(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_0),
    .D(GND_0),
    .Z(un1_main_basesoc_uart_rx_fifo_consume_c2_TMR_0)
  );
  defparam un1_main_basesoc_uart_rx_fifo_consume_ac0_1_TMR_0.INIT = "0x8080";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55826.8-55832.2" *)
  LUT4 un1_main_basesoc_uart_rx_fifo_consume_ac0_1_TMR_1 (
    .A(main_basesoc_uart_rx_fifo_consume_TMR_1[0]),
    .B(main_basesoc_uart_rx_fifo_consume_TMR_1[1]),
    .C(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_1),
    .D(GND_0),
    .Z(un1_main_basesoc_uart_rx_fifo_consume_c2_TMR_1)
  );
  defparam un1_main_basesoc_uart_rx_fifo_consume_ac0_1_TMR_1.INIT = "0x8080";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55826.8-55832.2" *)
  LUT4 un1_main_basesoc_uart_rx_fifo_consume_ac0_1_TMR_2 (
    .A(main_basesoc_uart_rx_fifo_consume_TMR_2[0]),
    .B(main_basesoc_uart_rx_fifo_consume_TMR_2[1]),
    .C(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_2),
    .D(GND_0),
    .Z(un1_main_basesoc_uart_rx_fifo_consume_c2_TMR_2)
  );
  defparam un1_main_basesoc_uart_rx_fifo_consume_ac0_1_TMR_2.INIT = "0x8080";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55853.8-55859.2" *)
  LUT4 un1_main_basesoc_uart_rx_fifo_consume_axbxc0_cZ_TMR_0 (
    .A(main_basesoc_uart_rx_fifo_consume_TMR_0[0]),
    .B(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_0),
    .C(GND_0),
    .D(GND_0),
    .Z(un1_main_basesoc_uart_rx_fifo_consume_axbxc0_TMR_0)
  );
  defparam un1_main_basesoc_uart_rx_fifo_consume_axbxc0_cZ_TMR_0.INIT = "0x6666";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55853.8-55859.2" *)
  LUT4 un1_main_basesoc_uart_rx_fifo_consume_axbxc0_cZ_TMR_1 (
    .A(main_basesoc_uart_rx_fifo_consume_TMR_1[0]),
    .B(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_1),
    .C(GND_0),
    .D(GND_0),
    .Z(un1_main_basesoc_uart_rx_fifo_consume_axbxc0_TMR_1)
  );
  defparam un1_main_basesoc_uart_rx_fifo_consume_axbxc0_cZ_TMR_1.INIT = "0x6666";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55853.8-55859.2" *)
  LUT4 un1_main_basesoc_uart_rx_fifo_consume_axbxc0_cZ_TMR_2 (
    .A(main_basesoc_uart_rx_fifo_consume_TMR_2[0]),
    .B(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_2),
    .C(GND_0),
    .D(GND_0),
    .Z(un1_main_basesoc_uart_rx_fifo_consume_axbxc0_TMR_2)
  );
  defparam un1_main_basesoc_uart_rx_fifo_consume_axbxc0_cZ_TMR_2.INIT = "0x6666";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55817.8-55823.2" *)
  LUT4 un1_main_basesoc_uart_rx_fifo_consume_axbxc1_cZ_TMR_0 (
    .A(main_basesoc_uart_rx_fifo_consume_TMR_0[0]),
    .B(main_basesoc_uart_rx_fifo_consume_TMR_0[1]),
    .C(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_0),
    .D(GND_0),
    .Z(un1_main_basesoc_uart_rx_fifo_consume_axbxc1_TMR_0)
  );
  defparam un1_main_basesoc_uart_rx_fifo_consume_axbxc1_cZ_TMR_0.INIT = "0x6C6C";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55817.8-55823.2" *)
  LUT4 un1_main_basesoc_uart_rx_fifo_consume_axbxc1_cZ_TMR_1 (
    .A(main_basesoc_uart_rx_fifo_consume_TMR_1[0]),
    .B(main_basesoc_uart_rx_fifo_consume_TMR_1[1]),
    .C(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_1),
    .D(GND_0),
    .Z(un1_main_basesoc_uart_rx_fifo_consume_axbxc1_TMR_1)
  );
  defparam un1_main_basesoc_uart_rx_fifo_consume_axbxc1_cZ_TMR_1.INIT = "0x6C6C";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55817.8-55823.2" *)
  LUT4 un1_main_basesoc_uart_rx_fifo_consume_axbxc1_cZ_TMR_2 (
    .A(main_basesoc_uart_rx_fifo_consume_TMR_2[0]),
    .B(main_basesoc_uart_rx_fifo_consume_TMR_2[1]),
    .C(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_2),
    .D(GND_0),
    .Z(un1_main_basesoc_uart_rx_fifo_consume_axbxc1_TMR_2)
  );
  defparam un1_main_basesoc_uart_rx_fifo_consume_axbxc1_cZ_TMR_2.INIT = "0x6C6C";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55665.8-55671.2" *)
  LUT4 un1_main_basesoc_uart_rx_fifo_consume_axbxc3_cZ_TMR_0 (
    .A(main_basesoc_uart_rx_fifo_consume_TMR_0[2]),
    .B(main_basesoc_uart_rx_fifo_consume_TMR_0[3]),
    .C(un1_main_basesoc_uart_rx_fifo_consume_c2_TMR_0),
    .D(GND_0),
    .Z(un1_main_basesoc_uart_rx_fifo_consume_axbxc3_TMR_0)
  );
  defparam un1_main_basesoc_uart_rx_fifo_consume_axbxc3_cZ_TMR_0.INIT = "0x6C6C";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55665.8-55671.2" *)
  LUT4 un1_main_basesoc_uart_rx_fifo_consume_axbxc3_cZ_TMR_1 (
    .A(main_basesoc_uart_rx_fifo_consume_TMR_1[2]),
    .B(main_basesoc_uart_rx_fifo_consume_TMR_1[3]),
    .C(un1_main_basesoc_uart_rx_fifo_consume_c2_TMR_1),
    .D(GND_0),
    .Z(un1_main_basesoc_uart_rx_fifo_consume_axbxc3_TMR_1)
  );
  defparam un1_main_basesoc_uart_rx_fifo_consume_axbxc3_cZ_TMR_1.INIT = "0x6C6C";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55665.8-55671.2" *)
  LUT4 un1_main_basesoc_uart_rx_fifo_consume_axbxc3_cZ_TMR_2 (
    .A(main_basesoc_uart_rx_fifo_consume_TMR_2[2]),
    .B(main_basesoc_uart_rx_fifo_consume_TMR_2[3]),
    .C(un1_main_basesoc_uart_rx_fifo_consume_c2_TMR_2),
    .D(GND_0),
    .Z(un1_main_basesoc_uart_rx_fifo_consume_axbxc3_TMR_2)
  );
  defparam un1_main_basesoc_uart_rx_fifo_consume_axbxc3_cZ_TMR_2.INIT = "0x6C6C";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56388.8-56401.2" *)
  CCU2 un1_main_basesoc_uart_rx_fifo_level0_cry_0_0_TMR_0 (
    .A0(VCC_TMR_0),
    .A1(un1_main_basesoc_uart_rx_fifo_level0_scalar_TMR_0),
    .B0(VCC_TMR_0),
    .B1(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_0),
    .C0(VCC_TMR_0),
    .C1(main_basesoc_uart_rx_fifo_wrport_we_TMR_0),
    .CIN(GND_0),
    .COUT(un1_main_basesoc_uart_rx_fifo_level0_cry_0_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un1_main_basesoc_uart_rx_fifo_level0_cry_0_0_S0_TMR_0),
    .S1(un1_main_basesoc_uart_rx_fifo_level0_cry_0_0_S1_TMR_0)
  );
  defparam un1_main_basesoc_uart_rx_fifo_level0_cry_0_0_TMR_0.INIT0 = "5033";
  defparam un1_main_basesoc_uart_rx_fifo_level0_cry_0_0_TMR_0.INIT1 = "96AA";
  defparam un1_main_basesoc_uart_rx_fifo_level0_cry_0_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56388.8-56401.2" *)
  CCU2 un1_main_basesoc_uart_rx_fifo_level0_cry_0_0_TMR_1 (
    .A0(VCC_TMR_1),
    .A1(un1_main_basesoc_uart_rx_fifo_level0_scalar_TMR_1),
    .B0(VCC_TMR_1),
    .B1(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_1),
    .C0(VCC_TMR_1),
    .C1(main_basesoc_uart_rx_fifo_wrport_we_TMR_1),
    .CIN(GND_0),
    .COUT(un1_main_basesoc_uart_rx_fifo_level0_cry_0_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un1_main_basesoc_uart_rx_fifo_level0_cry_0_0_S0_TMR_1),
    .S1(un1_main_basesoc_uart_rx_fifo_level0_cry_0_0_S1_TMR_1)
  );
  defparam un1_main_basesoc_uart_rx_fifo_level0_cry_0_0_TMR_1.INIT0 = "5033";
  defparam un1_main_basesoc_uart_rx_fifo_level0_cry_0_0_TMR_1.INIT1 = "96AA";
  defparam un1_main_basesoc_uart_rx_fifo_level0_cry_0_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56388.8-56401.2" *)
  CCU2 un1_main_basesoc_uart_rx_fifo_level0_cry_0_0_TMR_2 (
    .A0(VCC_TMR_2),
    .A1(un1_main_basesoc_uart_rx_fifo_level0_scalar_TMR_2),
    .B0(VCC_TMR_2),
    .B1(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_2),
    .C0(VCC_TMR_2),
    .C1(main_basesoc_uart_rx_fifo_wrport_we_TMR_2),
    .CIN(GND_0),
    .COUT(un1_main_basesoc_uart_rx_fifo_level0_cry_0_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un1_main_basesoc_uart_rx_fifo_level0_cry_0_0_S0_TMR_2),
    .S1(un1_main_basesoc_uart_rx_fifo_level0_cry_0_0_S1_TMR_2)
  );
  defparam un1_main_basesoc_uart_rx_fifo_level0_cry_0_0_TMR_2.INIT0 = "5033";
  defparam un1_main_basesoc_uart_rx_fifo_level0_cry_0_0_TMR_2.INIT1 = "96AA";
  defparam un1_main_basesoc_uart_rx_fifo_level0_cry_0_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56371.8-56384.2" *)
  CCU2 un1_main_basesoc_uart_rx_fifo_level0_cry_1_0_TMR_0 (
    .A0(un1_main_basesoc_uart_rx_fifo_level0_0_TMR_0[1]),
    .A1(un1_main_basesoc_uart_rx_fifo_level0_0_TMR_0[2]),
    .B0(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_0),
    .B1(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_0),
    .C0(main_basesoc_uart_rx_fifo_wrport_we_TMR_0),
    .C1(main_basesoc_uart_rx_fifo_wrport_we_TMR_0),
    .CIN(un1_main_basesoc_uart_rx_fifo_level0_cry_0_TMR_0),
    .COUT(un1_main_basesoc_uart_rx_fifo_level0_cry_2_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un1_main_basesoc_uart_rx_fifo_level0_TMR_0[1]),
    .S1(un1_main_basesoc_uart_rx_fifo_level0_TMR_0[2])
  );
  defparam un1_main_basesoc_uart_rx_fifo_level0_cry_1_0_TMR_0.INIT0 = "A6AA";
  defparam un1_main_basesoc_uart_rx_fifo_level0_cry_1_0_TMR_0.INIT1 = "A6AA";
  defparam un1_main_basesoc_uart_rx_fifo_level0_cry_1_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56371.8-56384.2" *)
  CCU2 un1_main_basesoc_uart_rx_fifo_level0_cry_1_0_TMR_1 (
    .A0(un1_main_basesoc_uart_rx_fifo_level0_0_TMR_1[1]),
    .A1(un1_main_basesoc_uart_rx_fifo_level0_0_TMR_1[2]),
    .B0(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_1),
    .B1(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_1),
    .C0(main_basesoc_uart_rx_fifo_wrport_we_TMR_1),
    .C1(main_basesoc_uart_rx_fifo_wrport_we_TMR_1),
    .CIN(un1_main_basesoc_uart_rx_fifo_level0_cry_0_TMR_1),
    .COUT(un1_main_basesoc_uart_rx_fifo_level0_cry_2_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un1_main_basesoc_uart_rx_fifo_level0_TMR_1[1]),
    .S1(un1_main_basesoc_uart_rx_fifo_level0_TMR_1[2])
  );
  defparam un1_main_basesoc_uart_rx_fifo_level0_cry_1_0_TMR_1.INIT0 = "A6AA";
  defparam un1_main_basesoc_uart_rx_fifo_level0_cry_1_0_TMR_1.INIT1 = "A6AA";
  defparam un1_main_basesoc_uart_rx_fifo_level0_cry_1_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56371.8-56384.2" *)
  CCU2 un1_main_basesoc_uart_rx_fifo_level0_cry_1_0_TMR_2 (
    .A0(un1_main_basesoc_uart_rx_fifo_level0_0_TMR_2[1]),
    .A1(un1_main_basesoc_uart_rx_fifo_level0_0_TMR_2[2]),
    .B0(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_2),
    .B1(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_2),
    .C0(main_basesoc_uart_rx_fifo_wrport_we_TMR_2),
    .C1(main_basesoc_uart_rx_fifo_wrport_we_TMR_2),
    .CIN(un1_main_basesoc_uart_rx_fifo_level0_cry_0_TMR_2),
    .COUT(un1_main_basesoc_uart_rx_fifo_level0_cry_2_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un1_main_basesoc_uart_rx_fifo_level0_TMR_2[1]),
    .S1(un1_main_basesoc_uart_rx_fifo_level0_TMR_2[2])
  );
  defparam un1_main_basesoc_uart_rx_fifo_level0_cry_1_0_TMR_2.INIT0 = "A6AA";
  defparam un1_main_basesoc_uart_rx_fifo_level0_cry_1_0_TMR_2.INIT1 = "A6AA";
  defparam un1_main_basesoc_uart_rx_fifo_level0_cry_1_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56353.8-56366.2" *)
  CCU2 un1_main_basesoc_uart_rx_fifo_level0_cry_3_0_TMR_0 (
    .A0(un1_main_basesoc_uart_rx_fifo_level0_0_TMR_0[3]),
    .A1(un1_main_basesoc_uart_rx_fifo_level0_0_TMR_0[4]),
    .B0(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_0),
    .B1(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_0),
    .C0(main_basesoc_uart_rx_fifo_wrport_we_TMR_0),
    .C1(main_basesoc_uart_rx_fifo_wrport_we_TMR_0),
    .CIN(un1_main_basesoc_uart_rx_fifo_level0_cry_2_TMR_0),
    .COUT(un1_main_basesoc_uart_rx_fifo_level0_cry_3_0_COUT_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un1_main_basesoc_uart_rx_fifo_level0_TMR_0[3]),
    .S1(un1_main_basesoc_uart_rx_fifo_level0_TMR_0[4])
  );
  defparam un1_main_basesoc_uart_rx_fifo_level0_cry_3_0_TMR_0.INIT0 = "A6AA";
  defparam un1_main_basesoc_uart_rx_fifo_level0_cry_3_0_TMR_0.INIT1 = "A6AA";
  defparam un1_main_basesoc_uart_rx_fifo_level0_cry_3_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56353.8-56366.2" *)
  CCU2 un1_main_basesoc_uart_rx_fifo_level0_cry_3_0_TMR_1 (
    .A0(un1_main_basesoc_uart_rx_fifo_level0_0_TMR_1[3]),
    .A1(un1_main_basesoc_uart_rx_fifo_level0_0_TMR_1[4]),
    .B0(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_1),
    .B1(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_1),
    .C0(main_basesoc_uart_rx_fifo_wrport_we_TMR_1),
    .C1(main_basesoc_uart_rx_fifo_wrport_we_TMR_1),
    .CIN(un1_main_basesoc_uart_rx_fifo_level0_cry_2_TMR_1),
    .COUT(un1_main_basesoc_uart_rx_fifo_level0_cry_3_0_COUT_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un1_main_basesoc_uart_rx_fifo_level0_TMR_1[3]),
    .S1(un1_main_basesoc_uart_rx_fifo_level0_TMR_1[4])
  );
  defparam un1_main_basesoc_uart_rx_fifo_level0_cry_3_0_TMR_1.INIT0 = "A6AA";
  defparam un1_main_basesoc_uart_rx_fifo_level0_cry_3_0_TMR_1.INIT1 = "A6AA";
  defparam un1_main_basesoc_uart_rx_fifo_level0_cry_3_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56353.8-56366.2" *)
  CCU2 un1_main_basesoc_uart_rx_fifo_level0_cry_3_0_TMR_2 (
    .A0(un1_main_basesoc_uart_rx_fifo_level0_0_TMR_2[3]),
    .A1(un1_main_basesoc_uart_rx_fifo_level0_0_TMR_2[4]),
    .B0(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_2),
    .B1(main_basesoc_uart_rx_fifo_syncfifo_re_TMR_2),
    .C0(main_basesoc_uart_rx_fifo_wrport_we_TMR_2),
    .C1(main_basesoc_uart_rx_fifo_wrport_we_TMR_2),
    .CIN(un1_main_basesoc_uart_rx_fifo_level0_cry_2_TMR_2),
    .COUT(un1_main_basesoc_uart_rx_fifo_level0_cry_3_0_COUT_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un1_main_basesoc_uart_rx_fifo_level0_TMR_2[3]),
    .S1(un1_main_basesoc_uart_rx_fifo_level0_TMR_2[4])
  );
  defparam un1_main_basesoc_uart_rx_fifo_level0_cry_3_0_TMR_2.INIT0 = "A6AA";
  defparam un1_main_basesoc_uart_rx_fifo_level0_cry_3_0_TMR_2.INIT1 = "A6AA";
  defparam un1_main_basesoc_uart_rx_fifo_level0_cry_3_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55791.8-55797.2" *)
  LUT4 un1_main_basesoc_uart_rx_fifo_produce_ac0_1_TMR_0 (
    .A(main_basesoc_uart_rx_fifo_produce_TMR_0[0]),
    .B(main_basesoc_uart_rx_fifo_produce_TMR_0[1]),
    .C(main_basesoc_uart_rx_fifo_wrport_we_TMR_0),
    .D(GND_0),
    .Z(un1_main_basesoc_uart_rx_fifo_produce_c2_TMR_0)
  );
  defparam un1_main_basesoc_uart_rx_fifo_produce_ac0_1_TMR_0.INIT = "0x8080";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55791.8-55797.2" *)
  LUT4 un1_main_basesoc_uart_rx_fifo_produce_ac0_1_TMR_1 (
    .A(main_basesoc_uart_rx_fifo_produce_TMR_1[0]),
    .B(main_basesoc_uart_rx_fifo_produce_TMR_1[1]),
    .C(main_basesoc_uart_rx_fifo_wrport_we_TMR_1),
    .D(GND_0),
    .Z(un1_main_basesoc_uart_rx_fifo_produce_c2_TMR_1)
  );
  defparam un1_main_basesoc_uart_rx_fifo_produce_ac0_1_TMR_1.INIT = "0x8080";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55791.8-55797.2" *)
  LUT4 un1_main_basesoc_uart_rx_fifo_produce_ac0_1_TMR_2 (
    .A(main_basesoc_uart_rx_fifo_produce_TMR_2[0]),
    .B(main_basesoc_uart_rx_fifo_produce_TMR_2[1]),
    .C(main_basesoc_uart_rx_fifo_wrport_we_TMR_2),
    .D(GND_0),
    .Z(un1_main_basesoc_uart_rx_fifo_produce_c2_TMR_2)
  );
  defparam un1_main_basesoc_uart_rx_fifo_produce_ac0_1_TMR_2.INIT = "0x8080";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55835.8-55841.2" *)
  LUT4 un1_main_basesoc_uart_rx_fifo_produce_axbxc0_cZ_TMR_0 (
    .A(main_basesoc_uart_rx_fifo_produce_TMR_0[0]),
    .B(main_basesoc_uart_rx_fifo_wrport_we_TMR_0),
    .C(GND_0),
    .D(GND_0),
    .Z(un1_main_basesoc_uart_rx_fifo_produce_axbxc0_TMR_0)
  );
  defparam un1_main_basesoc_uart_rx_fifo_produce_axbxc0_cZ_TMR_0.INIT = "0x6666";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55835.8-55841.2" *)
  LUT4 un1_main_basesoc_uart_rx_fifo_produce_axbxc0_cZ_TMR_1 (
    .A(main_basesoc_uart_rx_fifo_produce_TMR_1[0]),
    .B(main_basesoc_uart_rx_fifo_wrport_we_TMR_1),
    .C(GND_0),
    .D(GND_0),
    .Z(un1_main_basesoc_uart_rx_fifo_produce_axbxc0_TMR_1)
  );
  defparam un1_main_basesoc_uart_rx_fifo_produce_axbxc0_cZ_TMR_1.INIT = "0x6666";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55835.8-55841.2" *)
  LUT4 un1_main_basesoc_uart_rx_fifo_produce_axbxc0_cZ_TMR_2 (
    .A(main_basesoc_uart_rx_fifo_produce_TMR_2[0]),
    .B(main_basesoc_uart_rx_fifo_wrport_we_TMR_2),
    .C(GND_0),
    .D(GND_0),
    .Z(un1_main_basesoc_uart_rx_fifo_produce_axbxc0_TMR_2)
  );
  defparam un1_main_basesoc_uart_rx_fifo_produce_axbxc0_cZ_TMR_2.INIT = "0x6666";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55782.8-55788.2" *)
  LUT4 un1_main_basesoc_uart_rx_fifo_produce_axbxc1_cZ_TMR_0 (
    .A(main_basesoc_uart_rx_fifo_produce_TMR_0[0]),
    .B(main_basesoc_uart_rx_fifo_produce_TMR_0[1]),
    .C(main_basesoc_uart_rx_fifo_wrport_we_TMR_0),
    .D(GND_0),
    .Z(un1_main_basesoc_uart_rx_fifo_produce_axbxc1_TMR_0)
  );
  defparam un1_main_basesoc_uart_rx_fifo_produce_axbxc1_cZ_TMR_0.INIT = "0x6C6C";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55782.8-55788.2" *)
  LUT4 un1_main_basesoc_uart_rx_fifo_produce_axbxc1_cZ_TMR_1 (
    .A(main_basesoc_uart_rx_fifo_produce_TMR_1[0]),
    .B(main_basesoc_uart_rx_fifo_produce_TMR_1[1]),
    .C(main_basesoc_uart_rx_fifo_wrport_we_TMR_1),
    .D(GND_0),
    .Z(un1_main_basesoc_uart_rx_fifo_produce_axbxc1_TMR_1)
  );
  defparam un1_main_basesoc_uart_rx_fifo_produce_axbxc1_cZ_TMR_1.INIT = "0x6C6C";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55782.8-55788.2" *)
  LUT4 un1_main_basesoc_uart_rx_fifo_produce_axbxc1_cZ_TMR_2 (
    .A(main_basesoc_uart_rx_fifo_produce_TMR_2[0]),
    .B(main_basesoc_uart_rx_fifo_produce_TMR_2[1]),
    .C(main_basesoc_uart_rx_fifo_wrport_we_TMR_2),
    .D(GND_0),
    .Z(un1_main_basesoc_uart_rx_fifo_produce_axbxc1_TMR_2)
  );
  defparam un1_main_basesoc_uart_rx_fifo_produce_axbxc1_cZ_TMR_2.INIT = "0x6C6C";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55638.8-55644.2" *)
  LUT4 un1_main_basesoc_uart_rx_fifo_produce_axbxc3_cZ_TMR_0 (
    .A(main_basesoc_uart_rx_fifo_produce_TMR_0[2]),
    .B(main_basesoc_uart_rx_fifo_produce_TMR_0[3]),
    .C(un1_main_basesoc_uart_rx_fifo_produce_c2_TMR_0),
    .D(GND_0),
    .Z(un1_main_basesoc_uart_rx_fifo_produce_axbxc3_TMR_0)
  );
  defparam un1_main_basesoc_uart_rx_fifo_produce_axbxc3_cZ_TMR_0.INIT = "0x6C6C";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55638.8-55644.2" *)
  LUT4 un1_main_basesoc_uart_rx_fifo_produce_axbxc3_cZ_TMR_1 (
    .A(main_basesoc_uart_rx_fifo_produce_TMR_1[2]),
    .B(main_basesoc_uart_rx_fifo_produce_TMR_1[3]),
    .C(un1_main_basesoc_uart_rx_fifo_produce_c2_TMR_1),
    .D(GND_0),
    .Z(un1_main_basesoc_uart_rx_fifo_produce_axbxc3_TMR_1)
  );
  defparam un1_main_basesoc_uart_rx_fifo_produce_axbxc3_cZ_TMR_1.INIT = "0x6C6C";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55638.8-55644.2" *)
  LUT4 un1_main_basesoc_uart_rx_fifo_produce_axbxc3_cZ_TMR_2 (
    .A(main_basesoc_uart_rx_fifo_produce_TMR_2[2]),
    .B(main_basesoc_uart_rx_fifo_produce_TMR_2[3]),
    .C(un1_main_basesoc_uart_rx_fifo_produce_c2_TMR_2),
    .D(GND_0),
    .Z(un1_main_basesoc_uart_rx_fifo_produce_axbxc3_TMR_2)
  );
  defparam un1_main_basesoc_uart_rx_fifo_produce_axbxc3_cZ_TMR_2.INIT = "0x6C6C";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55683.8-55689.2" *)
  LUT4 un1_main_basesoc_uart_tx_fifo_consume_ac0_1_TMR_0 (
    .A(main_basesoc_uart_tx_fifo_consume_TMR_0[0]),
    .B(main_basesoc_uart_tx_fifo_consume_TMR_0[1]),
    .C(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_0),
    .D(GND_0),
    .Z(un1_main_basesoc_uart_tx_fifo_consume_c2_TMR_0)
  );
  defparam un1_main_basesoc_uart_tx_fifo_consume_ac0_1_TMR_0.INIT = "0x8080";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55683.8-55689.2" *)
  LUT4 un1_main_basesoc_uart_tx_fifo_consume_ac0_1_TMR_1 (
    .A(main_basesoc_uart_tx_fifo_consume_TMR_1[0]),
    .B(main_basesoc_uart_tx_fifo_consume_TMR_1[1]),
    .C(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_1),
    .D(GND_0),
    .Z(un1_main_basesoc_uart_tx_fifo_consume_c2_TMR_1)
  );
  defparam un1_main_basesoc_uart_tx_fifo_consume_ac0_1_TMR_1.INIT = "0x8080";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55683.8-55689.2" *)
  LUT4 un1_main_basesoc_uart_tx_fifo_consume_ac0_1_TMR_2 (
    .A(main_basesoc_uart_tx_fifo_consume_TMR_2[0]),
    .B(main_basesoc_uart_tx_fifo_consume_TMR_2[1]),
    .C(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_2),
    .D(GND_0),
    .Z(un1_main_basesoc_uart_tx_fifo_consume_c2_TMR_2)
  );
  defparam un1_main_basesoc_uart_tx_fifo_consume_ac0_1_TMR_2.INIT = "0x8080";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55773.8-55779.2" *)
  LUT4 un1_main_basesoc_uart_tx_fifo_consume_axbxc0_cZ_TMR_0 (
    .A(main_basesoc_uart_tx_fifo_consume_TMR_0[0]),
    .B(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_0),
    .C(GND_0),
    .D(GND_0),
    .Z(un1_main_basesoc_uart_tx_fifo_consume_axbxc0_TMR_0)
  );
  defparam un1_main_basesoc_uart_tx_fifo_consume_axbxc0_cZ_TMR_0.INIT = "0x6666";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55773.8-55779.2" *)
  LUT4 un1_main_basesoc_uart_tx_fifo_consume_axbxc0_cZ_TMR_1 (
    .A(main_basesoc_uart_tx_fifo_consume_TMR_1[0]),
    .B(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_1),
    .C(GND_0),
    .D(GND_0),
    .Z(un1_main_basesoc_uart_tx_fifo_consume_axbxc0_TMR_1)
  );
  defparam un1_main_basesoc_uart_tx_fifo_consume_axbxc0_cZ_TMR_1.INIT = "0x6666";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55773.8-55779.2" *)
  LUT4 un1_main_basesoc_uart_tx_fifo_consume_axbxc0_cZ_TMR_2 (
    .A(main_basesoc_uart_tx_fifo_consume_TMR_2[0]),
    .B(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_2),
    .C(GND_0),
    .D(GND_0),
    .Z(un1_main_basesoc_uart_tx_fifo_consume_axbxc0_TMR_2)
  );
  defparam un1_main_basesoc_uart_tx_fifo_consume_axbxc0_cZ_TMR_2.INIT = "0x6666";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55674.8-55680.2" *)
  LUT4 un1_main_basesoc_uart_tx_fifo_consume_axbxc1_cZ_TMR_0 (
    .A(main_basesoc_uart_tx_fifo_consume_TMR_0[0]),
    .B(main_basesoc_uart_tx_fifo_consume_TMR_0[1]),
    .C(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_0),
    .D(GND_0),
    .Z(un1_main_basesoc_uart_tx_fifo_consume_axbxc1_TMR_0)
  );
  defparam un1_main_basesoc_uart_tx_fifo_consume_axbxc1_cZ_TMR_0.INIT = "0x6C6C";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55674.8-55680.2" *)
  LUT4 un1_main_basesoc_uart_tx_fifo_consume_axbxc1_cZ_TMR_1 (
    .A(main_basesoc_uart_tx_fifo_consume_TMR_1[0]),
    .B(main_basesoc_uart_tx_fifo_consume_TMR_1[1]),
    .C(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_1),
    .D(GND_0),
    .Z(un1_main_basesoc_uart_tx_fifo_consume_axbxc1_TMR_1)
  );
  defparam un1_main_basesoc_uart_tx_fifo_consume_axbxc1_cZ_TMR_1.INIT = "0x6C6C";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55674.8-55680.2" *)
  LUT4 un1_main_basesoc_uart_tx_fifo_consume_axbxc1_cZ_TMR_2 (
    .A(main_basesoc_uart_tx_fifo_consume_TMR_2[0]),
    .B(main_basesoc_uart_tx_fifo_consume_TMR_2[1]),
    .C(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_2),
    .D(GND_0),
    .Z(un1_main_basesoc_uart_tx_fifo_consume_axbxc1_TMR_2)
  );
  defparam un1_main_basesoc_uart_tx_fifo_consume_axbxc1_cZ_TMR_2.INIT = "0x6C6C";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55613.8-55619.2" *)
  LUT4 un1_main_basesoc_uart_tx_fifo_consume_axbxc3_cZ_TMR_0 (
    .A(main_basesoc_uart_tx_fifo_consume_TMR_0[2]),
    .B(main_basesoc_uart_tx_fifo_consume_TMR_0[3]),
    .C(un1_main_basesoc_uart_tx_fifo_consume_c2_TMR_0),
    .D(GND_0),
    .Z(un1_main_basesoc_uart_tx_fifo_consume_axbxc3_TMR_0)
  );
  defparam un1_main_basesoc_uart_tx_fifo_consume_axbxc3_cZ_TMR_0.INIT = "0x6C6C";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55613.8-55619.2" *)
  LUT4 un1_main_basesoc_uart_tx_fifo_consume_axbxc3_cZ_TMR_1 (
    .A(main_basesoc_uart_tx_fifo_consume_TMR_1[2]),
    .B(main_basesoc_uart_tx_fifo_consume_TMR_1[3]),
    .C(un1_main_basesoc_uart_tx_fifo_consume_c2_TMR_1),
    .D(GND_0),
    .Z(un1_main_basesoc_uart_tx_fifo_consume_axbxc3_TMR_1)
  );
  defparam un1_main_basesoc_uart_tx_fifo_consume_axbxc3_cZ_TMR_1.INIT = "0x6C6C";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55613.8-55619.2" *)
  LUT4 un1_main_basesoc_uart_tx_fifo_consume_axbxc3_cZ_TMR_2 (
    .A(main_basesoc_uart_tx_fifo_consume_TMR_2[2]),
    .B(main_basesoc_uart_tx_fifo_consume_TMR_2[3]),
    .C(un1_main_basesoc_uart_tx_fifo_consume_c2_TMR_2),
    .D(GND_0),
    .Z(un1_main_basesoc_uart_tx_fifo_consume_axbxc3_TMR_2)
  );
  defparam un1_main_basesoc_uart_tx_fifo_consume_axbxc3_cZ_TMR_2.INIT = "0x6C6C";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56441.8-56454.2" *)
  CCU2 un1_main_basesoc_uart_tx_fifo_level0_cry_0_0_TMR_0 (
    .A0(VCC_TMR_0),
    .A1(un1_main_basesoc_uart_tx_fifo_level0_TMR_0[0]),
    .B0(VCC_TMR_0),
    .B1(un1_main_basesoc_uart_tx_fifo_level0_scalar_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(GND_0),
    .COUT(un1_main_basesoc_uart_tx_fifo_level0_cry_0_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un1_main_basesoc_uart_tx_fifo_level0_cry_0_0_S0_TMR_0),
    .S1(un1_main_basesoc_uart_tx_fifo_level0_cry_0_0_S1_TMR_0)
  );
  defparam un1_main_basesoc_uart_tx_fifo_level0_cry_0_0_TMR_0.INIT0 = "5033";
  defparam un1_main_basesoc_uart_tx_fifo_level0_cry_0_0_TMR_0.INIT1 = "A0CC";
  defparam un1_main_basesoc_uart_tx_fifo_level0_cry_0_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56441.8-56454.2" *)
  CCU2 un1_main_basesoc_uart_tx_fifo_level0_cry_0_0_TMR_1 (
    .A0(VCC_TMR_1),
    .A1(un1_main_basesoc_uart_tx_fifo_level0_TMR_1[0]),
    .B0(VCC_TMR_1),
    .B1(un1_main_basesoc_uart_tx_fifo_level0_scalar_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(GND_0),
    .COUT(un1_main_basesoc_uart_tx_fifo_level0_cry_0_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un1_main_basesoc_uart_tx_fifo_level0_cry_0_0_S0_TMR_1),
    .S1(un1_main_basesoc_uart_tx_fifo_level0_cry_0_0_S1_TMR_1)
  );
  defparam un1_main_basesoc_uart_tx_fifo_level0_cry_0_0_TMR_1.INIT0 = "5033";
  defparam un1_main_basesoc_uart_tx_fifo_level0_cry_0_0_TMR_1.INIT1 = "A0CC";
  defparam un1_main_basesoc_uart_tx_fifo_level0_cry_0_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56441.8-56454.2" *)
  CCU2 un1_main_basesoc_uart_tx_fifo_level0_cry_0_0_TMR_2 (
    .A0(VCC_TMR_2),
    .A1(un1_main_basesoc_uart_tx_fifo_level0_TMR_2[0]),
    .B0(VCC_TMR_2),
    .B1(un1_main_basesoc_uart_tx_fifo_level0_scalar_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(GND_0),
    .COUT(un1_main_basesoc_uart_tx_fifo_level0_cry_0_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un1_main_basesoc_uart_tx_fifo_level0_cry_0_0_S0_TMR_2),
    .S1(un1_main_basesoc_uart_tx_fifo_level0_cry_0_0_S1_TMR_2)
  );
  defparam un1_main_basesoc_uart_tx_fifo_level0_cry_0_0_TMR_2.INIT0 = "5033";
  defparam un1_main_basesoc_uart_tx_fifo_level0_cry_0_0_TMR_2.INIT1 = "A0CC";
  defparam un1_main_basesoc_uart_tx_fifo_level0_cry_0_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56424.8-56437.2" *)
  CCU2 un1_main_basesoc_uart_tx_fifo_level0_cry_1_0_TMR_0 (
    .A0(un1_main_basesoc_uart_tx_fifo_level0_0_TMR_0[1]),
    .A1(un1_main_basesoc_uart_tx_fifo_level0_0_TMR_0[2]),
    .B0(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_0),
    .B1(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_0),
    .C0(builder_csr_bankarray_interface0_bank_bus_dat_r8_6_RNIG6FO8_TMR_0),
    .C1(builder_csr_bankarray_interface0_bank_bus_dat_r8_6_RNIG6FO8_TMR_0),
    .CIN(un1_main_basesoc_uart_tx_fifo_level0_cry_0_TMR_0),
    .COUT(un1_main_basesoc_uart_tx_fifo_level0_cry_2_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un1_main_basesoc_uart_tx_fifo_level0_TMR_0[1]),
    .S1(un1_main_basesoc_uart_tx_fifo_level0_TMR_0[2])
  );
  defparam un1_main_basesoc_uart_tx_fifo_level0_cry_1_0_TMR_0.INIT0 = "A6AA";
  defparam un1_main_basesoc_uart_tx_fifo_level0_cry_1_0_TMR_0.INIT1 = "A6AA";
  defparam un1_main_basesoc_uart_tx_fifo_level0_cry_1_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56424.8-56437.2" *)
  CCU2 un1_main_basesoc_uart_tx_fifo_level0_cry_1_0_TMR_1 (
    .A0(un1_main_basesoc_uart_tx_fifo_level0_0_TMR_1[1]),
    .A1(un1_main_basesoc_uart_tx_fifo_level0_0_TMR_1[2]),
    .B0(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_1),
    .B1(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_1),
    .C0(builder_csr_bankarray_interface0_bank_bus_dat_r8_6_RNIG6FO8_TMR_1),
    .C1(builder_csr_bankarray_interface0_bank_bus_dat_r8_6_RNIG6FO8_TMR_1),
    .CIN(un1_main_basesoc_uart_tx_fifo_level0_cry_0_TMR_1),
    .COUT(un1_main_basesoc_uart_tx_fifo_level0_cry_2_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un1_main_basesoc_uart_tx_fifo_level0_TMR_1[1]),
    .S1(un1_main_basesoc_uart_tx_fifo_level0_TMR_1[2])
  );
  defparam un1_main_basesoc_uart_tx_fifo_level0_cry_1_0_TMR_1.INIT0 = "A6AA";
  defparam un1_main_basesoc_uart_tx_fifo_level0_cry_1_0_TMR_1.INIT1 = "A6AA";
  defparam un1_main_basesoc_uart_tx_fifo_level0_cry_1_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56424.8-56437.2" *)
  CCU2 un1_main_basesoc_uart_tx_fifo_level0_cry_1_0_TMR_2 (
    .A0(un1_main_basesoc_uart_tx_fifo_level0_0_TMR_2[1]),
    .A1(un1_main_basesoc_uart_tx_fifo_level0_0_TMR_2[2]),
    .B0(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_2),
    .B1(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_2),
    .C0(builder_csr_bankarray_interface0_bank_bus_dat_r8_6_RNIG6FO8_TMR_2),
    .C1(builder_csr_bankarray_interface0_bank_bus_dat_r8_6_RNIG6FO8_TMR_2),
    .CIN(un1_main_basesoc_uart_tx_fifo_level0_cry_0_TMR_2),
    .COUT(un1_main_basesoc_uart_tx_fifo_level0_cry_2_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un1_main_basesoc_uart_tx_fifo_level0_TMR_2[1]),
    .S1(un1_main_basesoc_uart_tx_fifo_level0_TMR_2[2])
  );
  defparam un1_main_basesoc_uart_tx_fifo_level0_cry_1_0_TMR_2.INIT0 = "A6AA";
  defparam un1_main_basesoc_uart_tx_fifo_level0_cry_1_0_TMR_2.INIT1 = "A6AA";
  defparam un1_main_basesoc_uart_tx_fifo_level0_cry_1_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56406.8-56419.2" *)
  CCU2 un1_main_basesoc_uart_tx_fifo_level0_cry_3_0_TMR_0 (
    .A0(un1_main_basesoc_uart_tx_fifo_level0_0_TMR_0[3]),
    .A1(un1_main_basesoc_uart_tx_fifo_level0_0_TMR_0[4]),
    .B0(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_0),
    .B1(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_0),
    .C0(builder_csr_bankarray_interface0_bank_bus_dat_r8_6_RNIG6FO8_TMR_0),
    .C1(builder_csr_bankarray_interface0_bank_bus_dat_r8_6_RNIG6FO8_TMR_0),
    .CIN(un1_main_basesoc_uart_tx_fifo_level0_cry_2_TMR_0),
    .COUT(un1_main_basesoc_uart_tx_fifo_level0_cry_3_0_COUT_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un1_main_basesoc_uart_tx_fifo_level0_TMR_0[3]),
    .S1(un1_main_basesoc_uart_tx_fifo_level0_TMR_0[4])
  );
  defparam un1_main_basesoc_uart_tx_fifo_level0_cry_3_0_TMR_0.INIT0 = "A6AA";
  defparam un1_main_basesoc_uart_tx_fifo_level0_cry_3_0_TMR_0.INIT1 = "A6AA";
  defparam un1_main_basesoc_uart_tx_fifo_level0_cry_3_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56406.8-56419.2" *)
  CCU2 un1_main_basesoc_uart_tx_fifo_level0_cry_3_0_TMR_1 (
    .A0(un1_main_basesoc_uart_tx_fifo_level0_0_TMR_1[3]),
    .A1(un1_main_basesoc_uart_tx_fifo_level0_0_TMR_1[4]),
    .B0(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_1),
    .B1(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_1),
    .C0(builder_csr_bankarray_interface0_bank_bus_dat_r8_6_RNIG6FO8_TMR_1),
    .C1(builder_csr_bankarray_interface0_bank_bus_dat_r8_6_RNIG6FO8_TMR_1),
    .CIN(un1_main_basesoc_uart_tx_fifo_level0_cry_2_TMR_1),
    .COUT(un1_main_basesoc_uart_tx_fifo_level0_cry_3_0_COUT_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un1_main_basesoc_uart_tx_fifo_level0_TMR_1[3]),
    .S1(un1_main_basesoc_uart_tx_fifo_level0_TMR_1[4])
  );
  defparam un1_main_basesoc_uart_tx_fifo_level0_cry_3_0_TMR_1.INIT0 = "A6AA";
  defparam un1_main_basesoc_uart_tx_fifo_level0_cry_3_0_TMR_1.INIT1 = "A6AA";
  defparam un1_main_basesoc_uart_tx_fifo_level0_cry_3_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56406.8-56419.2" *)
  CCU2 un1_main_basesoc_uart_tx_fifo_level0_cry_3_0_TMR_2 (
    .A0(un1_main_basesoc_uart_tx_fifo_level0_0_TMR_2[3]),
    .A1(un1_main_basesoc_uart_tx_fifo_level0_0_TMR_2[4]),
    .B0(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_2),
    .B1(main_basesoc_uart_tx_fifo_syncfifo_re_TMR_2),
    .C0(builder_csr_bankarray_interface0_bank_bus_dat_r8_6_RNIG6FO8_TMR_2),
    .C1(builder_csr_bankarray_interface0_bank_bus_dat_r8_6_RNIG6FO8_TMR_2),
    .CIN(un1_main_basesoc_uart_tx_fifo_level0_cry_2_TMR_2),
    .COUT(un1_main_basesoc_uart_tx_fifo_level0_cry_3_0_COUT_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un1_main_basesoc_uart_tx_fifo_level0_TMR_2[3]),
    .S1(un1_main_basesoc_uart_tx_fifo_level0_TMR_2[4])
  );
  defparam un1_main_basesoc_uart_tx_fifo_level0_cry_3_0_TMR_2.INIT0 = "A6AA";
  defparam un1_main_basesoc_uart_tx_fifo_level0_cry_3_0_TMR_2.INIT1 = "A6AA";
  defparam un1_main_basesoc_uart_tx_fifo_level0_cry_3_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55656.8-55662.2" *)
  LUT4 un1_main_basesoc_uart_tx_fifo_produce_ac0_0_cZ_TMR_0 (
    .A(N_167_TMR_0),
    .B(\VexRiscv.IBusCachedPlugin_cache.builder_slave_sel_r_r_0_a2_0_out_TMR_0 ),
    .C(\VexRiscv.main_m1_e_0_1_TMR_0 ),
    .D(main_basesoc_uart_tx_fifo_produce_TMR_0[0]),
    .Z(un1_main_basesoc_uart_tx_fifo_produce_ac0_0_TMR_0)
  );
  defparam un1_main_basesoc_uart_tx_fifo_produce_ac0_0_cZ_TMR_0.INIT = "0x8000";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55656.8-55662.2" *)
  LUT4 un1_main_basesoc_uart_tx_fifo_produce_ac0_0_cZ_TMR_1 (
    .A(N_167_TMR_1),
    .B(\VexRiscv.IBusCachedPlugin_cache.builder_slave_sel_r_r_0_a2_0_out_TMR_1 ),
    .C(\VexRiscv.main_m1_e_0_1_TMR_1 ),
    .D(main_basesoc_uart_tx_fifo_produce_TMR_1[0]),
    .Z(un1_main_basesoc_uart_tx_fifo_produce_ac0_0_TMR_1)
  );
  defparam un1_main_basesoc_uart_tx_fifo_produce_ac0_0_cZ_TMR_1.INIT = "0x8000";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55656.8-55662.2" *)
  LUT4 un1_main_basesoc_uart_tx_fifo_produce_ac0_0_cZ_TMR_2 (
    .A(N_167_TMR_2),
    .B(\VexRiscv.IBusCachedPlugin_cache.builder_slave_sel_r_r_0_a2_0_out_TMR_2 ),
    .C(\VexRiscv.main_m1_e_0_1_TMR_2 ),
    .D(main_basesoc_uart_tx_fifo_produce_TMR_2[0]),
    .Z(un1_main_basesoc_uart_tx_fifo_produce_ac0_0_TMR_2)
  );
  defparam un1_main_basesoc_uart_tx_fifo_produce_ac0_0_cZ_TMR_2.INIT = "0x8000";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56309.8-56315.2" *)
  LUT4 un1_main_basesoc_uart_tx_fifo_produce_axbxc0_cZ_TMR_0 (
    .A(\VexRiscv.main_m1_e_0_1_TMR_0 ),
    .B(builder_csr_bankarray_interface3_bank_bus_dat_r_0_sqmuxa_TMR_0),
    .C(main_basesoc_uart_tx_fifo_produce_TMR_0[0]),
    .D(GND_0),
    .Z(un1_main_basesoc_uart_tx_fifo_produce_axbxc0_TMR_0)
  );
  defparam un1_main_basesoc_uart_tx_fifo_produce_axbxc0_cZ_TMR_0.INIT = "0x7878";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56309.8-56315.2" *)
  LUT4 un1_main_basesoc_uart_tx_fifo_produce_axbxc0_cZ_TMR_1 (
    .A(\VexRiscv.main_m1_e_0_1_TMR_1 ),
    .B(builder_csr_bankarray_interface3_bank_bus_dat_r_0_sqmuxa_TMR_1),
    .C(main_basesoc_uart_tx_fifo_produce_TMR_1[0]),
    .D(GND_0),
    .Z(un1_main_basesoc_uart_tx_fifo_produce_axbxc0_TMR_1)
  );
  defparam un1_main_basesoc_uart_tx_fifo_produce_axbxc0_cZ_TMR_1.INIT = "0x7878";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56309.8-56315.2" *)
  LUT4 un1_main_basesoc_uart_tx_fifo_produce_axbxc0_cZ_TMR_2 (
    .A(\VexRiscv.main_m1_e_0_1_TMR_2 ),
    .B(builder_csr_bankarray_interface3_bank_bus_dat_r_0_sqmuxa_TMR_2),
    .C(main_basesoc_uart_tx_fifo_produce_TMR_2[0]),
    .D(GND_0),
    .Z(un1_main_basesoc_uart_tx_fifo_produce_axbxc0_TMR_2)
  );
  defparam un1_main_basesoc_uart_tx_fifo_produce_axbxc0_cZ_TMR_2.INIT = "0x7878";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55595.8-55601.2" *)
  LUT4 un1_main_basesoc_uart_tx_fifo_produce_axbxc1_cZ_TMR_0 (
    .A(builder_csr_bankarray_interface3_bank_bus_dat_r_0_sqmuxa_TMR_0),
    .B(main_basesoc_uart_tx_fifo_produce_TMR_0[1]),
    .C(un1_main_basesoc_uart_tx_fifo_produce_ac0_0_TMR_0),
    .D(GND_0),
    .Z(un1_main_basesoc_uart_tx_fifo_produce_axbxc1_TMR_0)
  );
  defparam un1_main_basesoc_uart_tx_fifo_produce_axbxc1_cZ_TMR_0.INIT = "0x6C6C";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55595.8-55601.2" *)
  LUT4 un1_main_basesoc_uart_tx_fifo_produce_axbxc1_cZ_TMR_1 (
    .A(builder_csr_bankarray_interface3_bank_bus_dat_r_0_sqmuxa_TMR_1),
    .B(main_basesoc_uart_tx_fifo_produce_TMR_1[1]),
    .C(un1_main_basesoc_uart_tx_fifo_produce_ac0_0_TMR_1),
    .D(GND_0),
    .Z(un1_main_basesoc_uart_tx_fifo_produce_axbxc1_TMR_1)
  );
  defparam un1_main_basesoc_uart_tx_fifo_produce_axbxc1_cZ_TMR_1.INIT = "0x6C6C";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55595.8-55601.2" *)
  LUT4 un1_main_basesoc_uart_tx_fifo_produce_axbxc1_cZ_TMR_2 (
    .A(builder_csr_bankarray_interface3_bank_bus_dat_r_0_sqmuxa_TMR_2),
    .B(main_basesoc_uart_tx_fifo_produce_TMR_2[1]),
    .C(un1_main_basesoc_uart_tx_fifo_produce_ac0_0_TMR_2),
    .D(GND_0),
    .Z(un1_main_basesoc_uart_tx_fifo_produce_axbxc1_TMR_2)
  );
  defparam un1_main_basesoc_uart_tx_fifo_produce_axbxc1_cZ_TMR_2.INIT = "0x6C6C";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55578.8-55584.2" *)
  LUT4 un1_main_basesoc_uart_tx_fifo_produce_axbxc2_cZ_TMR_0 (
    .A(builder_csr_bankarray_interface3_bank_bus_dat_r_0_sqmuxa_TMR_0),
    .B(main_basesoc_uart_tx_fifo_produce_TMR_0[1]),
    .C(main_basesoc_uart_tx_fifo_produce_TMR_0[2]),
    .D(un1_main_basesoc_uart_tx_fifo_produce_ac0_0_TMR_0),
    .Z(un1_main_basesoc_uart_tx_fifo_produce_axbxc2_TMR_0)
  );
  defparam un1_main_basesoc_uart_tx_fifo_produce_axbxc2_cZ_TMR_0.INIT = "0x78F0";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55578.8-55584.2" *)
  LUT4 un1_main_basesoc_uart_tx_fifo_produce_axbxc2_cZ_TMR_1 (
    .A(builder_csr_bankarray_interface3_bank_bus_dat_r_0_sqmuxa_TMR_1),
    .B(main_basesoc_uart_tx_fifo_produce_TMR_1[1]),
    .C(main_basesoc_uart_tx_fifo_produce_TMR_1[2]),
    .D(un1_main_basesoc_uart_tx_fifo_produce_ac0_0_TMR_1),
    .Z(un1_main_basesoc_uart_tx_fifo_produce_axbxc2_TMR_1)
  );
  defparam un1_main_basesoc_uart_tx_fifo_produce_axbxc2_cZ_TMR_1.INIT = "0x78F0";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55578.8-55584.2" *)
  LUT4 un1_main_basesoc_uart_tx_fifo_produce_axbxc2_cZ_TMR_2 (
    .A(builder_csr_bankarray_interface3_bank_bus_dat_r_0_sqmuxa_TMR_2),
    .B(main_basesoc_uart_tx_fifo_produce_TMR_2[1]),
    .C(main_basesoc_uart_tx_fifo_produce_TMR_2[2]),
    .D(un1_main_basesoc_uart_tx_fifo_produce_ac0_0_TMR_2),
    .Z(un1_main_basesoc_uart_tx_fifo_produce_axbxc2_TMR_2)
  );
  defparam un1_main_basesoc_uart_tx_fifo_produce_axbxc2_cZ_TMR_2.INIT = "0x78F0";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56264.8-56270.2" *)
  LUT4 un1_main_basesoc_uart_tx_fifo_produce_axbxc3_m6_e_0_cZ_TMR_0 (
    .A(main_basesoc_uart_tx_fifo_produce_TMR_0[1]),
    .B(main_basesoc_uart_tx_fifo_produce_TMR_0[2]),
    .C(GND_0),
    .D(GND_0),
    .Z(un1_main_basesoc_uart_tx_fifo_produce_axbxc3_m6_e_0_TMR_0)
  );
  defparam un1_main_basesoc_uart_tx_fifo_produce_axbxc3_m6_e_0_cZ_TMR_0.INIT = "0x8888";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56264.8-56270.2" *)
  LUT4 un1_main_basesoc_uart_tx_fifo_produce_axbxc3_m6_e_0_cZ_TMR_1 (
    .A(main_basesoc_uart_tx_fifo_produce_TMR_1[1]),
    .B(main_basesoc_uart_tx_fifo_produce_TMR_1[2]),
    .C(GND_0),
    .D(GND_0),
    .Z(un1_main_basesoc_uart_tx_fifo_produce_axbxc3_m6_e_0_TMR_1)
  );
  defparam un1_main_basesoc_uart_tx_fifo_produce_axbxc3_m6_e_0_cZ_TMR_1.INIT = "0x8888";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56264.8-56270.2" *)
  LUT4 un1_main_basesoc_uart_tx_fifo_produce_axbxc3_m6_e_0_cZ_TMR_2 (
    .A(main_basesoc_uart_tx_fifo_produce_TMR_2[1]),
    .B(main_basesoc_uart_tx_fifo_produce_TMR_2[2]),
    .C(GND_0),
    .D(GND_0),
    .Z(un1_main_basesoc_uart_tx_fifo_produce_axbxc3_m6_e_0_TMR_2)
  );
  defparam un1_main_basesoc_uart_tx_fifo_produce_axbxc3_m6_e_0_cZ_TMR_2.INIT = "0x8888";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55647.8-55653.2" *)
  LUT4 un1_main_basesoc_uart_tx_fifo_produce_axbxc3_m6_e_2_cZ_TMR_0 (
    .A(N_175_TMR_0),
    .B(\VexRiscv.builder_csr_bankarray_interface0_bank_bus_dat_r10_3_0_TMR_0 ),
    .C(main_basesoc_uart_tx_fifo_produce_TMR_0[0]),
    .D(un1_main_basesoc_uart_tx_fifo_produce_axbxc3_m6_e_0_TMR_0),
    .Z(un1_main_basesoc_uart_tx_fifo_produce_axbxc3_m6_e_2_TMR_0)
  );
  defparam un1_main_basesoc_uart_tx_fifo_produce_axbxc3_m6_e_2_cZ_TMR_0.INIT = "0xD000";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55647.8-55653.2" *)
  LUT4 un1_main_basesoc_uart_tx_fifo_produce_axbxc3_m6_e_2_cZ_TMR_1 (
    .A(N_175_TMR_1),
    .B(\VexRiscv.builder_csr_bankarray_interface0_bank_bus_dat_r10_3_0_TMR_1 ),
    .C(main_basesoc_uart_tx_fifo_produce_TMR_1[0]),
    .D(un1_main_basesoc_uart_tx_fifo_produce_axbxc3_m6_e_0_TMR_1),
    .Z(un1_main_basesoc_uart_tx_fifo_produce_axbxc3_m6_e_2_TMR_1)
  );
  defparam un1_main_basesoc_uart_tx_fifo_produce_axbxc3_m6_e_2_cZ_TMR_1.INIT = "0xD000";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55647.8-55653.2" *)
  LUT4 un1_main_basesoc_uart_tx_fifo_produce_axbxc3_m6_e_2_cZ_TMR_2 (
    .A(N_175_TMR_2),
    .B(\VexRiscv.builder_csr_bankarray_interface0_bank_bus_dat_r10_3_0_TMR_2 ),
    .C(main_basesoc_uart_tx_fifo_produce_TMR_2[0]),
    .D(un1_main_basesoc_uart_tx_fifo_produce_axbxc3_m6_e_0_TMR_2),
    .Z(un1_main_basesoc_uart_tx_fifo_produce_axbxc3_m6_e_2_TMR_2)
  );
  defparam un1_main_basesoc_uart_tx_fifo_produce_axbxc3_m6_e_2_cZ_TMR_2.INIT = "0xD000";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55604.8-55610.2" *)
  LUT4 un1_main_basesoc_uart_tx_fifo_produce_axbxc3_m6_e_TMR_0 (
    .A(\VexRiscv.builder_csr_bankarray_interface0_bank_bus_dat_r8_0_TMR_0 ),
    .B(un1_main_basesoc_uart_tx_fifo_produce_axbxc3_m6_e_2_TMR_0),
    .C(un1_main_basesoc_uart_tx_fifo_produce_axbxc3_m6_e_3_TMR_0),
    .D(GND_0),
    .Z(un1_main_basesoc_uart_tx_fifo_produce_axbxc3_N_13_mux_TMR_0)
  );
  defparam un1_main_basesoc_uart_tx_fifo_produce_axbxc3_m6_e_TMR_0.INIT = "0x8080";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55604.8-55610.2" *)
  LUT4 un1_main_basesoc_uart_tx_fifo_produce_axbxc3_m6_e_TMR_1 (
    .A(\VexRiscv.builder_csr_bankarray_interface0_bank_bus_dat_r8_0_TMR_1 ),
    .B(un1_main_basesoc_uart_tx_fifo_produce_axbxc3_m6_e_2_TMR_1),
    .C(un1_main_basesoc_uart_tx_fifo_produce_axbxc3_m6_e_3_TMR_1),
    .D(GND_0),
    .Z(un1_main_basesoc_uart_tx_fifo_produce_axbxc3_N_13_mux_TMR_1)
  );
  defparam un1_main_basesoc_uart_tx_fifo_produce_axbxc3_m6_e_TMR_1.INIT = "0x8080";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55604.8-55610.2" *)
  LUT4 un1_main_basesoc_uart_tx_fifo_produce_axbxc3_m6_e_TMR_2 (
    .A(\VexRiscv.builder_csr_bankarray_interface0_bank_bus_dat_r8_0_TMR_2 ),
    .B(un1_main_basesoc_uart_tx_fifo_produce_axbxc3_m6_e_2_TMR_2),
    .C(un1_main_basesoc_uart_tx_fifo_produce_axbxc3_m6_e_3_TMR_2),
    .D(GND_0),
    .Z(un1_main_basesoc_uart_tx_fifo_produce_axbxc3_N_13_mux_TMR_2)
  );
  defparam un1_main_basesoc_uart_tx_fifo_produce_axbxc3_m6_e_TMR_2.INIT = "0x8080";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56907.8-56920.2" *)
  CCU2 un1_main_crg_por_count_cry_0_0_TMR_0 (
    .A0(VCC_TMR_0),
    .A1(main_crg_por_count_TMR_0[0]),
    .B0(VCC_TMR_0),
    .B1(main_crg_por_done_13_TMR_0),
    .C0(VCC_TMR_0),
    .C1(main_crg_por_done_12_TMR_0),
    .CIN(GND_0),
    .COUT(un1_main_crg_por_count_cry_0_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un1_main_crg_por_count_cry_0_0_S0_TMR_0),
    .S1(un1_main_crg_por_count_cry_0_0_S1_TMR_0)
  );
  defparam un1_main_crg_por_count_cry_0_0_TMR_0.INIT0 = "5033";
  defparam un1_main_crg_por_count_cry_0_0_TMR_0.INIT1 = "95AA";
  defparam un1_main_crg_por_count_cry_0_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56907.8-56920.2" *)
  CCU2 un1_main_crg_por_count_cry_0_0_TMR_1 (
    .A0(VCC_TMR_1),
    .A1(main_crg_por_count_TMR_1[0]),
    .B0(VCC_TMR_1),
    .B1(main_crg_por_done_13_TMR_1),
    .C0(VCC_TMR_1),
    .C1(main_crg_por_done_12_TMR_1),
    .CIN(GND_0),
    .COUT(un1_main_crg_por_count_cry_0_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un1_main_crg_por_count_cry_0_0_S0_TMR_1),
    .S1(un1_main_crg_por_count_cry_0_0_S1_TMR_1)
  );
  defparam un1_main_crg_por_count_cry_0_0_TMR_1.INIT0 = "5033";
  defparam un1_main_crg_por_count_cry_0_0_TMR_1.INIT1 = "95AA";
  defparam un1_main_crg_por_count_cry_0_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56907.8-56920.2" *)
  CCU2 un1_main_crg_por_count_cry_0_0_TMR_2 (
    .A0(VCC_TMR_2),
    .A1(main_crg_por_count_TMR_2[0]),
    .B0(VCC_TMR_2),
    .B1(main_crg_por_done_13_TMR_2),
    .C0(VCC_TMR_2),
    .C1(main_crg_por_done_12_TMR_2),
    .CIN(GND_0),
    .COUT(un1_main_crg_por_count_cry_0_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un1_main_crg_por_count_cry_0_0_S0_TMR_2),
    .S1(un1_main_crg_por_count_cry_0_0_S1_TMR_2)
  );
  defparam un1_main_crg_por_count_cry_0_0_TMR_2.INIT0 = "5033";
  defparam un1_main_crg_por_count_cry_0_0_TMR_2.INIT1 = "95AA";
  defparam un1_main_crg_por_count_cry_0_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56800.8-56813.2" *)
  CCU2 un1_main_crg_por_count_cry_11_0_TMR_0 (
    .A0(main_crg_por_count_TMR_0[11]),
    .A1(main_crg_por_count_TMR_0[12]),
    .B0(main_crg_por_done_13_TMR_0),
    .B1(main_crg_por_done_13_TMR_0),
    .C0(main_crg_por_done_12_TMR_0),
    .C1(main_crg_por_done_12_TMR_0),
    .CIN(un1_main_crg_por_count_cry_10_TMR_0),
    .COUT(un1_main_crg_por_count_cry_12_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un1_main_crg_por_count_cry_11_0_S0_TMR_0),
    .S1(un1_main_crg_por_count_cry_11_0_S1_TMR_0)
  );
  defparam un1_main_crg_por_count_cry_11_0_TMR_0.INIT0 = "95AA";
  defparam un1_main_crg_por_count_cry_11_0_TMR_0.INIT1 = "95AA";
  defparam un1_main_crg_por_count_cry_11_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56800.8-56813.2" *)
  CCU2 un1_main_crg_por_count_cry_11_0_TMR_1 (
    .A0(main_crg_por_count_TMR_1[11]),
    .A1(main_crg_por_count_TMR_1[12]),
    .B0(main_crg_por_done_13_TMR_1),
    .B1(main_crg_por_done_13_TMR_1),
    .C0(main_crg_por_done_12_TMR_1),
    .C1(main_crg_por_done_12_TMR_1),
    .CIN(un1_main_crg_por_count_cry_10_TMR_1),
    .COUT(un1_main_crg_por_count_cry_12_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un1_main_crg_por_count_cry_11_0_S0_TMR_1),
    .S1(un1_main_crg_por_count_cry_11_0_S1_TMR_1)
  );
  defparam un1_main_crg_por_count_cry_11_0_TMR_1.INIT0 = "95AA";
  defparam un1_main_crg_por_count_cry_11_0_TMR_1.INIT1 = "95AA";
  defparam un1_main_crg_por_count_cry_11_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56800.8-56813.2" *)
  CCU2 un1_main_crg_por_count_cry_11_0_TMR_2 (
    .A0(main_crg_por_count_TMR_2[11]),
    .A1(main_crg_por_count_TMR_2[12]),
    .B0(main_crg_por_done_13_TMR_2),
    .B1(main_crg_por_done_13_TMR_2),
    .C0(main_crg_por_done_12_TMR_2),
    .C1(main_crg_por_done_12_TMR_2),
    .CIN(un1_main_crg_por_count_cry_10_TMR_2),
    .COUT(un1_main_crg_por_count_cry_12_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un1_main_crg_por_count_cry_11_0_S0_TMR_2),
    .S1(un1_main_crg_por_count_cry_11_0_S1_TMR_2)
  );
  defparam un1_main_crg_por_count_cry_11_0_TMR_2.INIT0 = "95AA";
  defparam un1_main_crg_por_count_cry_11_0_TMR_2.INIT1 = "95AA";
  defparam un1_main_crg_por_count_cry_11_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56782.8-56795.2" *)
  CCU2 un1_main_crg_por_count_cry_13_0_TMR_0 (
    .A0(main_crg_por_count_TMR_0[13]),
    .A1(main_crg_por_count_TMR_0[14]),
    .B0(main_crg_por_done_13_TMR_0),
    .B1(main_crg_por_done_13_TMR_0),
    .C0(main_crg_por_done_12_TMR_0),
    .C1(main_crg_por_done_12_TMR_0),
    .CIN(un1_main_crg_por_count_cry_12_TMR_0),
    .COUT(un1_main_crg_por_count_cry_14_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un1_main_crg_por_count_cry_13_0_S0_TMR_0),
    .S1(un1_main_crg_por_count_cry_13_0_S1_TMR_0)
  );
  defparam un1_main_crg_por_count_cry_13_0_TMR_0.INIT0 = "95AA";
  defparam un1_main_crg_por_count_cry_13_0_TMR_0.INIT1 = "95AA";
  defparam un1_main_crg_por_count_cry_13_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56782.8-56795.2" *)
  CCU2 un1_main_crg_por_count_cry_13_0_TMR_1 (
    .A0(main_crg_por_count_TMR_1[13]),
    .A1(main_crg_por_count_TMR_1[14]),
    .B0(main_crg_por_done_13_TMR_1),
    .B1(main_crg_por_done_13_TMR_1),
    .C0(main_crg_por_done_12_TMR_1),
    .C1(main_crg_por_done_12_TMR_1),
    .CIN(un1_main_crg_por_count_cry_12_TMR_1),
    .COUT(un1_main_crg_por_count_cry_14_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un1_main_crg_por_count_cry_13_0_S0_TMR_1),
    .S1(un1_main_crg_por_count_cry_13_0_S1_TMR_1)
  );
  defparam un1_main_crg_por_count_cry_13_0_TMR_1.INIT0 = "95AA";
  defparam un1_main_crg_por_count_cry_13_0_TMR_1.INIT1 = "95AA";
  defparam un1_main_crg_por_count_cry_13_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56782.8-56795.2" *)
  CCU2 un1_main_crg_por_count_cry_13_0_TMR_2 (
    .A0(main_crg_por_count_TMR_2[13]),
    .A1(main_crg_por_count_TMR_2[14]),
    .B0(main_crg_por_done_13_TMR_2),
    .B1(main_crg_por_done_13_TMR_2),
    .C0(main_crg_por_done_12_TMR_2),
    .C1(main_crg_por_done_12_TMR_2),
    .CIN(un1_main_crg_por_count_cry_12_TMR_2),
    .COUT(un1_main_crg_por_count_cry_14_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un1_main_crg_por_count_cry_13_0_S0_TMR_2),
    .S1(un1_main_crg_por_count_cry_13_0_S1_TMR_2)
  );
  defparam un1_main_crg_por_count_cry_13_0_TMR_2.INIT0 = "95AA";
  defparam un1_main_crg_por_count_cry_13_0_TMR_2.INIT1 = "95AA";
  defparam un1_main_crg_por_count_cry_13_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56890.8-56903.2" *)
  CCU2 un1_main_crg_por_count_cry_1_0_TMR_0 (
    .A0(main_crg_por_count_TMR_0[1]),
    .A1(main_crg_por_count_TMR_0[2]),
    .B0(main_crg_por_done_13_TMR_0),
    .B1(main_crg_por_done_13_TMR_0),
    .C0(main_crg_por_done_12_TMR_0),
    .C1(main_crg_por_done_12_TMR_0),
    .CIN(un1_main_crg_por_count_cry_0_TMR_0),
    .COUT(un1_main_crg_por_count_cry_2_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un1_main_crg_por_count_cry_1_0_S0_TMR_0),
    .S1(un1_main_crg_por_count_cry_1_0_S1_TMR_0)
  );
  defparam un1_main_crg_por_count_cry_1_0_TMR_0.INIT0 = "95AA";
  defparam un1_main_crg_por_count_cry_1_0_TMR_0.INIT1 = "95AA";
  defparam un1_main_crg_por_count_cry_1_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56890.8-56903.2" *)
  CCU2 un1_main_crg_por_count_cry_1_0_TMR_1 (
    .A0(main_crg_por_count_TMR_1[1]),
    .A1(main_crg_por_count_TMR_1[2]),
    .B0(main_crg_por_done_13_TMR_1),
    .B1(main_crg_por_done_13_TMR_1),
    .C0(main_crg_por_done_12_TMR_1),
    .C1(main_crg_por_done_12_TMR_1),
    .CIN(un1_main_crg_por_count_cry_0_TMR_1),
    .COUT(un1_main_crg_por_count_cry_2_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un1_main_crg_por_count_cry_1_0_S0_TMR_1),
    .S1(un1_main_crg_por_count_cry_1_0_S1_TMR_1)
  );
  defparam un1_main_crg_por_count_cry_1_0_TMR_1.INIT0 = "95AA";
  defparam un1_main_crg_por_count_cry_1_0_TMR_1.INIT1 = "95AA";
  defparam un1_main_crg_por_count_cry_1_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56890.8-56903.2" *)
  CCU2 un1_main_crg_por_count_cry_1_0_TMR_2 (
    .A0(main_crg_por_count_TMR_2[1]),
    .A1(main_crg_por_count_TMR_2[2]),
    .B0(main_crg_por_done_13_TMR_2),
    .B1(main_crg_por_done_13_TMR_2),
    .C0(main_crg_por_done_12_TMR_2),
    .C1(main_crg_por_done_12_TMR_2),
    .CIN(un1_main_crg_por_count_cry_0_TMR_2),
    .COUT(un1_main_crg_por_count_cry_2_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un1_main_crg_por_count_cry_1_0_S0_TMR_2),
    .S1(un1_main_crg_por_count_cry_1_0_S1_TMR_2)
  );
  defparam un1_main_crg_por_count_cry_1_0_TMR_2.INIT0 = "95AA";
  defparam un1_main_crg_por_count_cry_1_0_TMR_2.INIT1 = "95AA";
  defparam un1_main_crg_por_count_cry_1_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56872.8-56885.2" *)
  CCU2 un1_main_crg_por_count_cry_3_0_TMR_0 (
    .A0(main_crg_por_count_TMR_0[3]),
    .A1(main_crg_por_count_TMR_0[4]),
    .B0(main_crg_por_done_13_TMR_0),
    .B1(main_crg_por_done_13_TMR_0),
    .C0(main_crg_por_done_12_TMR_0),
    .C1(main_crg_por_done_12_TMR_0),
    .CIN(un1_main_crg_por_count_cry_2_TMR_0),
    .COUT(un1_main_crg_por_count_cry_4_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un1_main_crg_por_count_cry_3_0_S0_TMR_0),
    .S1(un1_main_crg_por_count_cry_3_0_S1_TMR_0)
  );
  defparam un1_main_crg_por_count_cry_3_0_TMR_0.INIT0 = "95AA";
  defparam un1_main_crg_por_count_cry_3_0_TMR_0.INIT1 = "95AA";
  defparam un1_main_crg_por_count_cry_3_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56872.8-56885.2" *)
  CCU2 un1_main_crg_por_count_cry_3_0_TMR_1 (
    .A0(main_crg_por_count_TMR_1[3]),
    .A1(main_crg_por_count_TMR_1[4]),
    .B0(main_crg_por_done_13_TMR_1),
    .B1(main_crg_por_done_13_TMR_1),
    .C0(main_crg_por_done_12_TMR_1),
    .C1(main_crg_por_done_12_TMR_1),
    .CIN(un1_main_crg_por_count_cry_2_TMR_1),
    .COUT(un1_main_crg_por_count_cry_4_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un1_main_crg_por_count_cry_3_0_S0_TMR_1),
    .S1(un1_main_crg_por_count_cry_3_0_S1_TMR_1)
  );
  defparam un1_main_crg_por_count_cry_3_0_TMR_1.INIT0 = "95AA";
  defparam un1_main_crg_por_count_cry_3_0_TMR_1.INIT1 = "95AA";
  defparam un1_main_crg_por_count_cry_3_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56872.8-56885.2" *)
  CCU2 un1_main_crg_por_count_cry_3_0_TMR_2 (
    .A0(main_crg_por_count_TMR_2[3]),
    .A1(main_crg_por_count_TMR_2[4]),
    .B0(main_crg_por_done_13_TMR_2),
    .B1(main_crg_por_done_13_TMR_2),
    .C0(main_crg_por_done_12_TMR_2),
    .C1(main_crg_por_done_12_TMR_2),
    .CIN(un1_main_crg_por_count_cry_2_TMR_2),
    .COUT(un1_main_crg_por_count_cry_4_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un1_main_crg_por_count_cry_3_0_S0_TMR_2),
    .S1(un1_main_crg_por_count_cry_3_0_S1_TMR_2)
  );
  defparam un1_main_crg_por_count_cry_3_0_TMR_2.INIT0 = "95AA";
  defparam un1_main_crg_por_count_cry_3_0_TMR_2.INIT1 = "95AA";
  defparam un1_main_crg_por_count_cry_3_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56854.8-56867.2" *)
  CCU2 un1_main_crg_por_count_cry_5_0_TMR_0 (
    .A0(main_crg_por_count_TMR_0[5]),
    .A1(main_crg_por_count_TMR_0[6]),
    .B0(main_crg_por_done_13_TMR_0),
    .B1(main_crg_por_done_13_TMR_0),
    .C0(main_crg_por_done_12_TMR_0),
    .C1(main_crg_por_done_12_TMR_0),
    .CIN(un1_main_crg_por_count_cry_4_TMR_0),
    .COUT(un1_main_crg_por_count_cry_6_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un1_main_crg_por_count_cry_5_0_S0_TMR_0),
    .S1(un1_main_crg_por_count_cry_5_0_S1_TMR_0)
  );
  defparam un1_main_crg_por_count_cry_5_0_TMR_0.INIT0 = "95AA";
  defparam un1_main_crg_por_count_cry_5_0_TMR_0.INIT1 = "95AA";
  defparam un1_main_crg_por_count_cry_5_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56854.8-56867.2" *)
  CCU2 un1_main_crg_por_count_cry_5_0_TMR_1 (
    .A0(main_crg_por_count_TMR_1[5]),
    .A1(main_crg_por_count_TMR_1[6]),
    .B0(main_crg_por_done_13_TMR_1),
    .B1(main_crg_por_done_13_TMR_1),
    .C0(main_crg_por_done_12_TMR_1),
    .C1(main_crg_por_done_12_TMR_1),
    .CIN(un1_main_crg_por_count_cry_4_TMR_1),
    .COUT(un1_main_crg_por_count_cry_6_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un1_main_crg_por_count_cry_5_0_S0_TMR_1),
    .S1(un1_main_crg_por_count_cry_5_0_S1_TMR_1)
  );
  defparam un1_main_crg_por_count_cry_5_0_TMR_1.INIT0 = "95AA";
  defparam un1_main_crg_por_count_cry_5_0_TMR_1.INIT1 = "95AA";
  defparam un1_main_crg_por_count_cry_5_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56854.8-56867.2" *)
  CCU2 un1_main_crg_por_count_cry_5_0_TMR_2 (
    .A0(main_crg_por_count_TMR_2[5]),
    .A1(main_crg_por_count_TMR_2[6]),
    .B0(main_crg_por_done_13_TMR_2),
    .B1(main_crg_por_done_13_TMR_2),
    .C0(main_crg_por_done_12_TMR_2),
    .C1(main_crg_por_done_12_TMR_2),
    .CIN(un1_main_crg_por_count_cry_4_TMR_2),
    .COUT(un1_main_crg_por_count_cry_6_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un1_main_crg_por_count_cry_5_0_S0_TMR_2),
    .S1(un1_main_crg_por_count_cry_5_0_S1_TMR_2)
  );
  defparam un1_main_crg_por_count_cry_5_0_TMR_2.INIT0 = "95AA";
  defparam un1_main_crg_por_count_cry_5_0_TMR_2.INIT1 = "95AA";
  defparam un1_main_crg_por_count_cry_5_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56836.8-56849.2" *)
  CCU2 un1_main_crg_por_count_cry_7_0_TMR_0 (
    .A0(main_crg_por_count_TMR_0[7]),
    .A1(main_crg_por_count_TMR_0[8]),
    .B0(main_crg_por_done_13_TMR_0),
    .B1(main_crg_por_done_13_TMR_0),
    .C0(main_crg_por_done_12_TMR_0),
    .C1(main_crg_por_done_12_TMR_0),
    .CIN(un1_main_crg_por_count_cry_6_TMR_0),
    .COUT(un1_main_crg_por_count_cry_8_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un1_main_crg_por_count_cry_7_0_S0_TMR_0),
    .S1(un1_main_crg_por_count_cry_7_0_S1_TMR_0)
  );
  defparam un1_main_crg_por_count_cry_7_0_TMR_0.INIT0 = "95AA";
  defparam un1_main_crg_por_count_cry_7_0_TMR_0.INIT1 = "95AA";
  defparam un1_main_crg_por_count_cry_7_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56836.8-56849.2" *)
  CCU2 un1_main_crg_por_count_cry_7_0_TMR_1 (
    .A0(main_crg_por_count_TMR_1[7]),
    .A1(main_crg_por_count_TMR_1[8]),
    .B0(main_crg_por_done_13_TMR_1),
    .B1(main_crg_por_done_13_TMR_1),
    .C0(main_crg_por_done_12_TMR_1),
    .C1(main_crg_por_done_12_TMR_1),
    .CIN(un1_main_crg_por_count_cry_6_TMR_1),
    .COUT(un1_main_crg_por_count_cry_8_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un1_main_crg_por_count_cry_7_0_S0_TMR_1),
    .S1(un1_main_crg_por_count_cry_7_0_S1_TMR_1)
  );
  defparam un1_main_crg_por_count_cry_7_0_TMR_1.INIT0 = "95AA";
  defparam un1_main_crg_por_count_cry_7_0_TMR_1.INIT1 = "95AA";
  defparam un1_main_crg_por_count_cry_7_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56836.8-56849.2" *)
  CCU2 un1_main_crg_por_count_cry_7_0_TMR_2 (
    .A0(main_crg_por_count_TMR_2[7]),
    .A1(main_crg_por_count_TMR_2[8]),
    .B0(main_crg_por_done_13_TMR_2),
    .B1(main_crg_por_done_13_TMR_2),
    .C0(main_crg_por_done_12_TMR_2),
    .C1(main_crg_por_done_12_TMR_2),
    .CIN(un1_main_crg_por_count_cry_6_TMR_2),
    .COUT(un1_main_crg_por_count_cry_8_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un1_main_crg_por_count_cry_7_0_S0_TMR_2),
    .S1(un1_main_crg_por_count_cry_7_0_S1_TMR_2)
  );
  defparam un1_main_crg_por_count_cry_7_0_TMR_2.INIT0 = "95AA";
  defparam un1_main_crg_por_count_cry_7_0_TMR_2.INIT1 = "95AA";
  defparam un1_main_crg_por_count_cry_7_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56818.8-56831.2" *)
  CCU2 un1_main_crg_por_count_cry_9_0_TMR_0 (
    .A0(main_crg_por_count_TMR_0[9]),
    .A1(main_crg_por_count_TMR_0[10]),
    .B0(main_crg_por_done_13_TMR_0),
    .B1(main_crg_por_done_13_TMR_0),
    .C0(main_crg_por_done_12_TMR_0),
    .C1(main_crg_por_done_12_TMR_0),
    .CIN(un1_main_crg_por_count_cry_8_TMR_0),
    .COUT(un1_main_crg_por_count_cry_10_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un1_main_crg_por_count_cry_9_0_S0_TMR_0),
    .S1(un1_main_crg_por_count_cry_9_0_S1_TMR_0)
  );
  defparam un1_main_crg_por_count_cry_9_0_TMR_0.INIT0 = "95AA";
  defparam un1_main_crg_por_count_cry_9_0_TMR_0.INIT1 = "95AA";
  defparam un1_main_crg_por_count_cry_9_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56818.8-56831.2" *)
  CCU2 un1_main_crg_por_count_cry_9_0_TMR_1 (
    .A0(main_crg_por_count_TMR_1[9]),
    .A1(main_crg_por_count_TMR_1[10]),
    .B0(main_crg_por_done_13_TMR_1),
    .B1(main_crg_por_done_13_TMR_1),
    .C0(main_crg_por_done_12_TMR_1),
    .C1(main_crg_por_done_12_TMR_1),
    .CIN(un1_main_crg_por_count_cry_8_TMR_1),
    .COUT(un1_main_crg_por_count_cry_10_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un1_main_crg_por_count_cry_9_0_S0_TMR_1),
    .S1(un1_main_crg_por_count_cry_9_0_S1_TMR_1)
  );
  defparam un1_main_crg_por_count_cry_9_0_TMR_1.INIT0 = "95AA";
  defparam un1_main_crg_por_count_cry_9_0_TMR_1.INIT1 = "95AA";
  defparam un1_main_crg_por_count_cry_9_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56818.8-56831.2" *)
  CCU2 un1_main_crg_por_count_cry_9_0_TMR_2 (
    .A0(main_crg_por_count_TMR_2[9]),
    .A1(main_crg_por_count_TMR_2[10]),
    .B0(main_crg_por_done_13_TMR_2),
    .B1(main_crg_por_done_13_TMR_2),
    .C0(main_crg_por_done_12_TMR_2),
    .C1(main_crg_por_done_12_TMR_2),
    .CIN(un1_main_crg_por_count_cry_8_TMR_2),
    .COUT(un1_main_crg_por_count_cry_10_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un1_main_crg_por_count_cry_9_0_S0_TMR_2),
    .S1(un1_main_crg_por_count_cry_9_0_S1_TMR_2)
  );
  defparam un1_main_crg_por_count_cry_9_0_TMR_2.INIT0 = "95AA";
  defparam un1_main_crg_por_count_cry_9_0_TMR_2.INIT1 = "95AA";
  defparam un1_main_crg_por_count_cry_9_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56764.8-56777.2" *)
  CCU2 un1_main_crg_por_count_s_15_0_TMR_0 (
    .A0(main_crg_por_count_TMR_0[15]),
    .A1(VCC_TMR_0),
    .B0(main_crg_por_done_13_TMR_0),
    .B1(VCC_TMR_0),
    .C0(main_crg_por_done_12_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(un1_main_crg_por_count_cry_14_TMR_0),
    .COUT(un1_main_crg_por_count_s_15_0_COUT_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un1_main_crg_por_count_s_15_0_S0_TMR_0),
    .S1(un1_main_crg_por_count_s_15_0_S1_TMR_0)
  );
  defparam un1_main_crg_por_count_s_15_0_TMR_0.INIT0 = "95AA";
  defparam un1_main_crg_por_count_s_15_0_TMR_0.INIT1 = "5033";
  defparam un1_main_crg_por_count_s_15_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56764.8-56777.2" *)
  CCU2 un1_main_crg_por_count_s_15_0_TMR_1 (
    .A0(main_crg_por_count_TMR_1[15]),
    .A1(VCC_TMR_1),
    .B0(main_crg_por_done_13_TMR_1),
    .B1(VCC_TMR_1),
    .C0(main_crg_por_done_12_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(un1_main_crg_por_count_cry_14_TMR_1),
    .COUT(un1_main_crg_por_count_s_15_0_COUT_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un1_main_crg_por_count_s_15_0_S0_TMR_1),
    .S1(un1_main_crg_por_count_s_15_0_S1_TMR_1)
  );
  defparam un1_main_crg_por_count_s_15_0_TMR_1.INIT0 = "95AA";
  defparam un1_main_crg_por_count_s_15_0_TMR_1.INIT1 = "5033";
  defparam un1_main_crg_por_count_s_15_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56764.8-56777.2" *)
  CCU2 un1_main_crg_por_count_s_15_0_TMR_2 (
    .A0(main_crg_por_count_TMR_2[15]),
    .A1(VCC_TMR_2),
    .B0(main_crg_por_done_13_TMR_2),
    .B1(VCC_TMR_2),
    .C0(main_crg_por_done_12_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(un1_main_crg_por_count_cry_14_TMR_2),
    .COUT(un1_main_crg_por_count_s_15_0_COUT_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un1_main_crg_por_count_s_15_0_S0_TMR_2),
    .S1(un1_main_crg_por_count_s_15_0_S1_TMR_2)
  );
  defparam un1_main_crg_por_count_s_15_0_TMR_2.INIT0 = "95AA";
  defparam un1_main_crg_por_count_s_15_0_TMR_2.INIT1 = "5033";
  defparam un1_main_crg_por_count_s_15_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55844.8-55850.2" *)
  LUT4 un2_main_crg_por_done_1_cZ_TMR_0 (
    .A(main_crg_locked),
    .B(main_crg_por_done_12_TMR_0),
    .C(main_crg_por_done_13_TMR_0),
    .D(GND_0),
    .Z(un2_main_crg_por_done_1_TMR_0)
  );
  defparam un2_main_crg_por_done_1_cZ_TMR_0.INIT = "0x7F7F";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55844.8-55850.2" *)
  LUT4 un2_main_crg_por_done_1_cZ_TMR_1 (
    .A(main_crg_locked),
    .B(main_crg_por_done_12_TMR_1),
    .C(main_crg_por_done_13_TMR_1),
    .D(GND_0),
    .Z(un2_main_crg_por_done_1_TMR_1)
  );
  defparam un2_main_crg_por_done_1_cZ_TMR_1.INIT = "0x7F7F";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55844.8-55850.2" *)
  LUT4 un2_main_crg_por_done_1_cZ_TMR_2 (
    .A(main_crg_locked),
    .B(main_crg_por_done_12_TMR_2),
    .C(main_crg_por_done_13_TMR_2),
    .D(GND_0),
    .Z(un2_main_crg_por_done_1_TMR_2)
  );
  defparam un2_main_crg_por_done_1_cZ_TMR_2.INIT = "0x7F7F";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57212.8-57225.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_0_0_TMR_0 (
    .A0(VCC_TMR_0),
    .A1(dsp_join_kb_27_TMR_0[0]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(GND_0),
    .COUT(un5_main_basesoc_rx_phase_cry_0_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un5_main_basesoc_rx_phase_cry_0_0_S0_TMR_0),
    .S1(un5_main_basesoc_rx_phase_cry_0_0_S1_TMR_0)
  );
  defparam un5_main_basesoc_rx_phase_cry_0_0_TMR_0.INIT0 = "5033";
  defparam un5_main_basesoc_rx_phase_cry_0_0_TMR_0.INIT1 = "50AA";
  defparam un5_main_basesoc_rx_phase_cry_0_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57212.8-57225.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_0_0_TMR_1 (
    .A0(VCC_TMR_1),
    .A1(dsp_join_kb_27_TMR_1[0]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(GND_0),
    .COUT(un5_main_basesoc_rx_phase_cry_0_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un5_main_basesoc_rx_phase_cry_0_0_S0_TMR_1),
    .S1(un5_main_basesoc_rx_phase_cry_0_0_S1_TMR_1)
  );
  defparam un5_main_basesoc_rx_phase_cry_0_0_TMR_1.INIT0 = "5033";
  defparam un5_main_basesoc_rx_phase_cry_0_0_TMR_1.INIT1 = "50AA";
  defparam un5_main_basesoc_rx_phase_cry_0_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57212.8-57225.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_0_0_TMR_2 (
    .A0(VCC_TMR_2),
    .A1(dsp_join_kb_27_TMR_2[0]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(GND_0),
    .COUT(un5_main_basesoc_rx_phase_cry_0_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un5_main_basesoc_rx_phase_cry_0_0_S0_TMR_2),
    .S1(un5_main_basesoc_rx_phase_cry_0_0_S1_TMR_2)
  );
  defparam un5_main_basesoc_rx_phase_cry_0_0_TMR_2.INIT0 = "5033";
  defparam un5_main_basesoc_rx_phase_cry_0_0_TMR_2.INIT1 = "50AA";
  defparam un5_main_basesoc_rx_phase_cry_0_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57105.8-57118.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_11_0_TMR_0 (
    .A0(dsp_join_kb_27_TMR_0[11]),
    .A1(dsp_join_kb_27_TMR_0[12]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(un5_main_basesoc_rx_phase_cry_10_TMR_0),
    .COUT(un5_main_basesoc_rx_phase_cry_12_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(N_413_TMR_0),
    .S1(N_414_TMR_0)
  );
  defparam un5_main_basesoc_rx_phase_cry_11_0_TMR_0.INIT0 = "50AA";
  defparam un5_main_basesoc_rx_phase_cry_11_0_TMR_0.INIT1 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_11_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57105.8-57118.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_11_0_TMR_1 (
    .A0(dsp_join_kb_27_TMR_1[11]),
    .A1(dsp_join_kb_27_TMR_1[12]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(un5_main_basesoc_rx_phase_cry_10_TMR_1),
    .COUT(un5_main_basesoc_rx_phase_cry_12_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(N_413_TMR_1),
    .S1(N_414_TMR_1)
  );
  defparam un5_main_basesoc_rx_phase_cry_11_0_TMR_1.INIT0 = "50AA";
  defparam un5_main_basesoc_rx_phase_cry_11_0_TMR_1.INIT1 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_11_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57105.8-57118.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_11_0_TMR_2 (
    .A0(dsp_join_kb_27_TMR_2[11]),
    .A1(dsp_join_kb_27_TMR_2[12]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(un5_main_basesoc_rx_phase_cry_10_TMR_2),
    .COUT(un5_main_basesoc_rx_phase_cry_12_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(N_413_TMR_2),
    .S1(N_414_TMR_2)
  );
  defparam un5_main_basesoc_rx_phase_cry_11_0_TMR_2.INIT0 = "50AA";
  defparam un5_main_basesoc_rx_phase_cry_11_0_TMR_2.INIT1 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_11_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57087.8-57100.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_13_0_TMR_0 (
    .A0(dsp_join_kb_27_TMR_0[13]),
    .A1(dsp_join_kb_27_TMR_0[14]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(un5_main_basesoc_rx_phase_cry_12_TMR_0),
    .COUT(un5_main_basesoc_rx_phase_cry_14_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(N_415_TMR_0),
    .S1(N_416_TMR_0)
  );
  defparam un5_main_basesoc_rx_phase_cry_13_0_TMR_0.INIT0 = "50AA";
  defparam un5_main_basesoc_rx_phase_cry_13_0_TMR_0.INIT1 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_13_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57087.8-57100.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_13_0_TMR_1 (
    .A0(dsp_join_kb_27_TMR_1[13]),
    .A1(dsp_join_kb_27_TMR_1[14]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(un5_main_basesoc_rx_phase_cry_12_TMR_1),
    .COUT(un5_main_basesoc_rx_phase_cry_14_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(N_415_TMR_1),
    .S1(N_416_TMR_1)
  );
  defparam un5_main_basesoc_rx_phase_cry_13_0_TMR_1.INIT0 = "50AA";
  defparam un5_main_basesoc_rx_phase_cry_13_0_TMR_1.INIT1 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_13_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57087.8-57100.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_13_0_TMR_2 (
    .A0(dsp_join_kb_27_TMR_2[13]),
    .A1(dsp_join_kb_27_TMR_2[14]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(un5_main_basesoc_rx_phase_cry_12_TMR_2),
    .COUT(un5_main_basesoc_rx_phase_cry_14_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(N_415_TMR_2),
    .S1(N_416_TMR_2)
  );
  defparam un5_main_basesoc_rx_phase_cry_13_0_TMR_2.INIT0 = "50AA";
  defparam un5_main_basesoc_rx_phase_cry_13_0_TMR_2.INIT1 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_13_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57069.8-57082.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_15_0_TMR_0 (
    .A0(dsp_join_kb_27_TMR_0[15]),
    .A1(dsp_join_kb_27_TMR_0[16]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(un5_main_basesoc_rx_phase_cry_14_TMR_0),
    .COUT(un5_main_basesoc_rx_phase_cry_16_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(N_417_TMR_0),
    .S1(un5_main_basesoc_rx_phase_cry_15_0_S1_TMR_0)
  );
  defparam un5_main_basesoc_rx_phase_cry_15_0_TMR_0.INIT0 = "50AA";
  defparam un5_main_basesoc_rx_phase_cry_15_0_TMR_0.INIT1 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_15_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57069.8-57082.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_15_0_TMR_1 (
    .A0(dsp_join_kb_27_TMR_1[15]),
    .A1(dsp_join_kb_27_TMR_1[16]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(un5_main_basesoc_rx_phase_cry_14_TMR_1),
    .COUT(un5_main_basesoc_rx_phase_cry_16_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(N_417_TMR_1),
    .S1(un5_main_basesoc_rx_phase_cry_15_0_S1_TMR_1)
  );
  defparam un5_main_basesoc_rx_phase_cry_15_0_TMR_1.INIT0 = "50AA";
  defparam un5_main_basesoc_rx_phase_cry_15_0_TMR_1.INIT1 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_15_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57069.8-57082.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_15_0_TMR_2 (
    .A0(dsp_join_kb_27_TMR_2[15]),
    .A1(dsp_join_kb_27_TMR_2[16]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(un5_main_basesoc_rx_phase_cry_14_TMR_2),
    .COUT(un5_main_basesoc_rx_phase_cry_16_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(N_417_TMR_2),
    .S1(un5_main_basesoc_rx_phase_cry_15_0_S1_TMR_2)
  );
  defparam un5_main_basesoc_rx_phase_cry_15_0_TMR_2.INIT0 = "50AA";
  defparam un5_main_basesoc_rx_phase_cry_15_0_TMR_2.INIT1 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_15_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57051.8-57064.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_17_0_TMR_0 (
    .A0(dsp_join_kb_27_TMR_0[17]),
    .A1(dsp_join_kb_27_TMR_0[18]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(un5_main_basesoc_rx_phase_cry_16_TMR_0),
    .COUT(un5_main_basesoc_rx_phase_cry_18_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(N_419_TMR_0),
    .S1(N_420_TMR_0)
  );
  defparam un5_main_basesoc_rx_phase_cry_17_0_TMR_0.INIT0 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_17_0_TMR_0.INIT1 = "50AA";
  defparam un5_main_basesoc_rx_phase_cry_17_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57051.8-57064.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_17_0_TMR_1 (
    .A0(dsp_join_kb_27_TMR_1[17]),
    .A1(dsp_join_kb_27_TMR_1[18]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(un5_main_basesoc_rx_phase_cry_16_TMR_1),
    .COUT(un5_main_basesoc_rx_phase_cry_18_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(N_419_TMR_1),
    .S1(N_420_TMR_1)
  );
  defparam un5_main_basesoc_rx_phase_cry_17_0_TMR_1.INIT0 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_17_0_TMR_1.INIT1 = "50AA";
  defparam un5_main_basesoc_rx_phase_cry_17_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57051.8-57064.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_17_0_TMR_2 (
    .A0(dsp_join_kb_27_TMR_2[17]),
    .A1(dsp_join_kb_27_TMR_2[18]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(un5_main_basesoc_rx_phase_cry_16_TMR_2),
    .COUT(un5_main_basesoc_rx_phase_cry_18_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(N_419_TMR_2),
    .S1(N_420_TMR_2)
  );
  defparam un5_main_basesoc_rx_phase_cry_17_0_TMR_2.INIT0 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_17_0_TMR_2.INIT1 = "50AA";
  defparam un5_main_basesoc_rx_phase_cry_17_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57033.8-57046.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_19_0_TMR_0 (
    .A0(dsp_join_kb_27_TMR_0[19]),
    .A1(dsp_join_kb_27_TMR_0[20]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(un5_main_basesoc_rx_phase_cry_18_TMR_0),
    .COUT(un5_main_basesoc_rx_phase_cry_20_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un5_main_basesoc_rx_phase_cry_19_0_S0_TMR_0),
    .S1(un5_main_basesoc_rx_phase_cry_19_0_S1_TMR_0)
  );
  defparam un5_main_basesoc_rx_phase_cry_19_0_TMR_0.INIT0 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_19_0_TMR_0.INIT1 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_19_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57033.8-57046.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_19_0_TMR_1 (
    .A0(dsp_join_kb_27_TMR_1[19]),
    .A1(dsp_join_kb_27_TMR_1[20]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(un5_main_basesoc_rx_phase_cry_18_TMR_1),
    .COUT(un5_main_basesoc_rx_phase_cry_20_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un5_main_basesoc_rx_phase_cry_19_0_S0_TMR_1),
    .S1(un5_main_basesoc_rx_phase_cry_19_0_S1_TMR_1)
  );
  defparam un5_main_basesoc_rx_phase_cry_19_0_TMR_1.INIT0 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_19_0_TMR_1.INIT1 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_19_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57033.8-57046.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_19_0_TMR_2 (
    .A0(dsp_join_kb_27_TMR_2[19]),
    .A1(dsp_join_kb_27_TMR_2[20]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(un5_main_basesoc_rx_phase_cry_18_TMR_2),
    .COUT(un5_main_basesoc_rx_phase_cry_20_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un5_main_basesoc_rx_phase_cry_19_0_S0_TMR_2),
    .S1(un5_main_basesoc_rx_phase_cry_19_0_S1_TMR_2)
  );
  defparam un5_main_basesoc_rx_phase_cry_19_0_TMR_2.INIT0 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_19_0_TMR_2.INIT1 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_19_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57195.8-57208.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_1_0_TMR_0 (
    .A0(dsp_join_kb_27_TMR_0[1]),
    .A1(dsp_join_kb_27_TMR_0[2]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(un5_main_basesoc_rx_phase_cry_0_TMR_0),
    .COUT(un5_main_basesoc_rx_phase_cry_2_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(N_403_TMR_0),
    .S1(N_404_TMR_0)
  );
  defparam un5_main_basesoc_rx_phase_cry_1_0_TMR_0.INIT0 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_1_0_TMR_0.INIT1 = "50AA";
  defparam un5_main_basesoc_rx_phase_cry_1_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57195.8-57208.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_1_0_TMR_1 (
    .A0(dsp_join_kb_27_TMR_1[1]),
    .A1(dsp_join_kb_27_TMR_1[2]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(un5_main_basesoc_rx_phase_cry_0_TMR_1),
    .COUT(un5_main_basesoc_rx_phase_cry_2_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(N_403_TMR_1),
    .S1(N_404_TMR_1)
  );
  defparam un5_main_basesoc_rx_phase_cry_1_0_TMR_1.INIT0 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_1_0_TMR_1.INIT1 = "50AA";
  defparam un5_main_basesoc_rx_phase_cry_1_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57195.8-57208.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_1_0_TMR_2 (
    .A0(dsp_join_kb_27_TMR_2[1]),
    .A1(dsp_join_kb_27_TMR_2[2]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(un5_main_basesoc_rx_phase_cry_0_TMR_2),
    .COUT(un5_main_basesoc_rx_phase_cry_2_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(N_403_TMR_2),
    .S1(N_404_TMR_2)
  );
  defparam un5_main_basesoc_rx_phase_cry_1_0_TMR_2.INIT0 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_1_0_TMR_2.INIT1 = "50AA";
  defparam un5_main_basesoc_rx_phase_cry_1_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57015.8-57028.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_21_0_TMR_0 (
    .A0(dsp_join_kb_27_TMR_0[21]),
    .A1(dsp_join_kb_27_TMR_0[22]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(un5_main_basesoc_rx_phase_cry_20_TMR_0),
    .COUT(un5_main_basesoc_rx_phase_cry_22_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(N_423_TMR_0),
    .S1(N_424_TMR_0)
  );
  defparam un5_main_basesoc_rx_phase_cry_21_0_TMR_0.INIT0 = "50AA";
  defparam un5_main_basesoc_rx_phase_cry_21_0_TMR_0.INIT1 = "50AA";
  defparam un5_main_basesoc_rx_phase_cry_21_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57015.8-57028.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_21_0_TMR_1 (
    .A0(dsp_join_kb_27_TMR_1[21]),
    .A1(dsp_join_kb_27_TMR_1[22]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(un5_main_basesoc_rx_phase_cry_20_TMR_1),
    .COUT(un5_main_basesoc_rx_phase_cry_22_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(N_423_TMR_1),
    .S1(N_424_TMR_1)
  );
  defparam un5_main_basesoc_rx_phase_cry_21_0_TMR_1.INIT0 = "50AA";
  defparam un5_main_basesoc_rx_phase_cry_21_0_TMR_1.INIT1 = "50AA";
  defparam un5_main_basesoc_rx_phase_cry_21_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57015.8-57028.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_21_0_TMR_2 (
    .A0(dsp_join_kb_27_TMR_2[21]),
    .A1(dsp_join_kb_27_TMR_2[22]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(un5_main_basesoc_rx_phase_cry_20_TMR_2),
    .COUT(un5_main_basesoc_rx_phase_cry_22_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(N_423_TMR_2),
    .S1(N_424_TMR_2)
  );
  defparam un5_main_basesoc_rx_phase_cry_21_0_TMR_2.INIT0 = "50AA";
  defparam un5_main_basesoc_rx_phase_cry_21_0_TMR_2.INIT1 = "50AA";
  defparam un5_main_basesoc_rx_phase_cry_21_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56997.8-57010.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_23_0_TMR_0 (
    .A0(dsp_join_kb_27_TMR_0[23]),
    .A1(dsp_join_kb_27_TMR_0[24]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(un5_main_basesoc_rx_phase_cry_22_TMR_0),
    .COUT(un5_main_basesoc_rx_phase_cry_24_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(N_425_TMR_0),
    .S1(un5_main_basesoc_rx_phase_cry_23_0_S1_TMR_0)
  );
  defparam un5_main_basesoc_rx_phase_cry_23_0_TMR_0.INIT0 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_23_0_TMR_0.INIT1 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_23_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56997.8-57010.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_23_0_TMR_1 (
    .A0(dsp_join_kb_27_TMR_1[23]),
    .A1(dsp_join_kb_27_TMR_1[24]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(un5_main_basesoc_rx_phase_cry_22_TMR_1),
    .COUT(un5_main_basesoc_rx_phase_cry_24_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(N_425_TMR_1),
    .S1(un5_main_basesoc_rx_phase_cry_23_0_S1_TMR_1)
  );
  defparam un5_main_basesoc_rx_phase_cry_23_0_TMR_1.INIT0 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_23_0_TMR_1.INIT1 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_23_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56997.8-57010.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_23_0_TMR_2 (
    .A0(dsp_join_kb_27_TMR_2[23]),
    .A1(dsp_join_kb_27_TMR_2[24]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(un5_main_basesoc_rx_phase_cry_22_TMR_2),
    .COUT(un5_main_basesoc_rx_phase_cry_24_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(N_425_TMR_2),
    .S1(un5_main_basesoc_rx_phase_cry_23_0_S1_TMR_2)
  );
  defparam un5_main_basesoc_rx_phase_cry_23_0_TMR_2.INIT0 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_23_0_TMR_2.INIT1 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_23_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56979.8-56992.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_25_0_TMR_0 (
    .A0(dsp_join_kb_27_TMR_0[25]),
    .A1(dsp_join_kb_27_TMR_0[26]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(un5_main_basesoc_rx_phase_cry_24_TMR_0),
    .COUT(un5_main_basesoc_rx_phase_cry_26_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(N_427_TMR_0),
    .S1(N_428_TMR_0)
  );
  defparam un5_main_basesoc_rx_phase_cry_25_0_TMR_0.INIT0 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_25_0_TMR_0.INIT1 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_25_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56979.8-56992.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_25_0_TMR_1 (
    .A0(dsp_join_kb_27_TMR_1[25]),
    .A1(dsp_join_kb_27_TMR_1[26]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(un5_main_basesoc_rx_phase_cry_24_TMR_1),
    .COUT(un5_main_basesoc_rx_phase_cry_26_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(N_427_TMR_1),
    .S1(N_428_TMR_1)
  );
  defparam un5_main_basesoc_rx_phase_cry_25_0_TMR_1.INIT0 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_25_0_TMR_1.INIT1 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_25_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56979.8-56992.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_25_0_TMR_2 (
    .A0(dsp_join_kb_27_TMR_2[25]),
    .A1(dsp_join_kb_27_TMR_2[26]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(un5_main_basesoc_rx_phase_cry_24_TMR_2),
    .COUT(un5_main_basesoc_rx_phase_cry_26_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(N_427_TMR_2),
    .S1(N_428_TMR_2)
  );
  defparam un5_main_basesoc_rx_phase_cry_25_0_TMR_2.INIT0 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_25_0_TMR_2.INIT1 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_25_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56961.8-56974.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_27_0_TMR_0 (
    .A0(dsp_join_kb_27_TMR_0[27]),
    .A1(dsp_join_kb_27_TMR_0[28]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(un5_main_basesoc_rx_phase_cry_26_TMR_0),
    .COUT(un5_main_basesoc_rx_phase_cry_28_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(N_429_TMR_0),
    .S1(N_430_TMR_0)
  );
  defparam un5_main_basesoc_rx_phase_cry_27_0_TMR_0.INIT0 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_27_0_TMR_0.INIT1 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_27_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56961.8-56974.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_27_0_TMR_1 (
    .A0(dsp_join_kb_27_TMR_1[27]),
    .A1(dsp_join_kb_27_TMR_1[28]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(un5_main_basesoc_rx_phase_cry_26_TMR_1),
    .COUT(un5_main_basesoc_rx_phase_cry_28_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(N_429_TMR_1),
    .S1(N_430_TMR_1)
  );
  defparam un5_main_basesoc_rx_phase_cry_27_0_TMR_1.INIT0 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_27_0_TMR_1.INIT1 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_27_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56961.8-56974.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_27_0_TMR_2 (
    .A0(dsp_join_kb_27_TMR_2[27]),
    .A1(dsp_join_kb_27_TMR_2[28]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(un5_main_basesoc_rx_phase_cry_26_TMR_2),
    .COUT(un5_main_basesoc_rx_phase_cry_28_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(N_429_TMR_2),
    .S1(N_430_TMR_2)
  );
  defparam un5_main_basesoc_rx_phase_cry_27_0_TMR_2.INIT0 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_27_0_TMR_2.INIT1 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_27_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56943.8-56956.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_29_0_TMR_0 (
    .A0(dsp_join_kb_27_TMR_0[29]),
    .A1(dsp_join_kb_27_TMR_0[30]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(un5_main_basesoc_rx_phase_cry_28_TMR_0),
    .COUT(un5_main_basesoc_rx_phase_cry_30_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un5_main_basesoc_rx_phase_cry_29_0_S0_TMR_0),
    .S1(un5_main_basesoc_rx_phase_cry_29_0_S1_TMR_0)
  );
  defparam un5_main_basesoc_rx_phase_cry_29_0_TMR_0.INIT0 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_29_0_TMR_0.INIT1 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_29_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56943.8-56956.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_29_0_TMR_1 (
    .A0(dsp_join_kb_27_TMR_1[29]),
    .A1(dsp_join_kb_27_TMR_1[30]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(un5_main_basesoc_rx_phase_cry_28_TMR_1),
    .COUT(un5_main_basesoc_rx_phase_cry_30_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un5_main_basesoc_rx_phase_cry_29_0_S0_TMR_1),
    .S1(un5_main_basesoc_rx_phase_cry_29_0_S1_TMR_1)
  );
  defparam un5_main_basesoc_rx_phase_cry_29_0_TMR_1.INIT0 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_29_0_TMR_1.INIT1 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_29_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56943.8-56956.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_29_0_TMR_2 (
    .A0(dsp_join_kb_27_TMR_2[29]),
    .A1(dsp_join_kb_27_TMR_2[30]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(un5_main_basesoc_rx_phase_cry_28_TMR_2),
    .COUT(un5_main_basesoc_rx_phase_cry_30_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un5_main_basesoc_rx_phase_cry_29_0_S0_TMR_2),
    .S1(un5_main_basesoc_rx_phase_cry_29_0_S1_TMR_2)
  );
  defparam un5_main_basesoc_rx_phase_cry_29_0_TMR_2.INIT0 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_29_0_TMR_2.INIT1 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_29_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56925.8-56938.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_31_0_TMR_0 (
    .A0(dsp_join_kb_27_TMR_0[31]),
    .A1(VCC_TMR_0),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(un5_main_basesoc_rx_phase_cry_30_TMR_0),
    .COUT(un5_main_basesoc_rx_phase_cry_31_0_COUT_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un5_main_basesoc_rx_phase_cry_31_0_S0_TMR_0),
    .S1(un5_main_basesoc_rx_phase_cry_31_TMR_0)
  );
  defparam un5_main_basesoc_rx_phase_cry_31_0_TMR_0.INIT0 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_31_0_TMR_0.INIT1 = "5033";
  defparam un5_main_basesoc_rx_phase_cry_31_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56925.8-56938.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_31_0_TMR_1 (
    .A0(dsp_join_kb_27_TMR_1[31]),
    .A1(VCC_TMR_1),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(un5_main_basesoc_rx_phase_cry_30_TMR_1),
    .COUT(un5_main_basesoc_rx_phase_cry_31_0_COUT_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un5_main_basesoc_rx_phase_cry_31_0_S0_TMR_1),
    .S1(un5_main_basesoc_rx_phase_cry_31_TMR_1)
  );
  defparam un5_main_basesoc_rx_phase_cry_31_0_TMR_1.INIT0 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_31_0_TMR_1.INIT1 = "5033";
  defparam un5_main_basesoc_rx_phase_cry_31_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:56925.8-56938.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_31_0_TMR_2 (
    .A0(dsp_join_kb_27_TMR_2[31]),
    .A1(VCC_TMR_2),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(un5_main_basesoc_rx_phase_cry_30_TMR_2),
    .COUT(un5_main_basesoc_rx_phase_cry_31_0_COUT_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un5_main_basesoc_rx_phase_cry_31_0_S0_TMR_2),
    .S1(un5_main_basesoc_rx_phase_cry_31_TMR_2)
  );
  defparam un5_main_basesoc_rx_phase_cry_31_0_TMR_2.INIT0 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_31_0_TMR_2.INIT1 = "5033";
  defparam un5_main_basesoc_rx_phase_cry_31_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57177.8-57190.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_3_0_TMR_0 (
    .A0(dsp_join_kb_27_TMR_0[3]),
    .A1(dsp_join_kb_27_TMR_0[4]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(un5_main_basesoc_rx_phase_cry_2_TMR_0),
    .COUT(un5_main_basesoc_rx_phase_cry_4_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(N_405_TMR_0),
    .S1(N_406_TMR_0)
  );
  defparam un5_main_basesoc_rx_phase_cry_3_0_TMR_0.INIT0 = "50AA";
  defparam un5_main_basesoc_rx_phase_cry_3_0_TMR_0.INIT1 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_3_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57177.8-57190.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_3_0_TMR_1 (
    .A0(dsp_join_kb_27_TMR_1[3]),
    .A1(dsp_join_kb_27_TMR_1[4]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(un5_main_basesoc_rx_phase_cry_2_TMR_1),
    .COUT(un5_main_basesoc_rx_phase_cry_4_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(N_405_TMR_1),
    .S1(N_406_TMR_1)
  );
  defparam un5_main_basesoc_rx_phase_cry_3_0_TMR_1.INIT0 = "50AA";
  defparam un5_main_basesoc_rx_phase_cry_3_0_TMR_1.INIT1 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_3_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57177.8-57190.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_3_0_TMR_2 (
    .A0(dsp_join_kb_27_TMR_2[3]),
    .A1(dsp_join_kb_27_TMR_2[4]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(un5_main_basesoc_rx_phase_cry_2_TMR_2),
    .COUT(un5_main_basesoc_rx_phase_cry_4_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(N_405_TMR_2),
    .S1(N_406_TMR_2)
  );
  defparam un5_main_basesoc_rx_phase_cry_3_0_TMR_2.INIT0 = "50AA";
  defparam un5_main_basesoc_rx_phase_cry_3_0_TMR_2.INIT1 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_3_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57159.8-57172.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_5_0_TMR_0 (
    .A0(dsp_join_kb_27_TMR_0[5]),
    .A1(dsp_join_kb_27_TMR_0[6]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(un5_main_basesoc_rx_phase_cry_4_TMR_0),
    .COUT(un5_main_basesoc_rx_phase_cry_6_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(N_407_TMR_0),
    .S1(N_408_TMR_0)
  );
  defparam un5_main_basesoc_rx_phase_cry_5_0_TMR_0.INIT0 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_5_0_TMR_0.INIT1 = "50AA";
  defparam un5_main_basesoc_rx_phase_cry_5_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57159.8-57172.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_5_0_TMR_1 (
    .A0(dsp_join_kb_27_TMR_1[5]),
    .A1(dsp_join_kb_27_TMR_1[6]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(un5_main_basesoc_rx_phase_cry_4_TMR_1),
    .COUT(un5_main_basesoc_rx_phase_cry_6_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(N_407_TMR_1),
    .S1(N_408_TMR_1)
  );
  defparam un5_main_basesoc_rx_phase_cry_5_0_TMR_1.INIT0 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_5_0_TMR_1.INIT1 = "50AA";
  defparam un5_main_basesoc_rx_phase_cry_5_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57159.8-57172.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_5_0_TMR_2 (
    .A0(dsp_join_kb_27_TMR_2[5]),
    .A1(dsp_join_kb_27_TMR_2[6]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(un5_main_basesoc_rx_phase_cry_4_TMR_2),
    .COUT(un5_main_basesoc_rx_phase_cry_6_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(N_407_TMR_2),
    .S1(N_408_TMR_2)
  );
  defparam un5_main_basesoc_rx_phase_cry_5_0_TMR_2.INIT0 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_5_0_TMR_2.INIT1 = "50AA";
  defparam un5_main_basesoc_rx_phase_cry_5_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57141.8-57154.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_7_0_TMR_0 (
    .A0(dsp_join_kb_27_TMR_0[7]),
    .A1(dsp_join_kb_27_TMR_0[8]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(un5_main_basesoc_rx_phase_cry_6_TMR_0),
    .COUT(un5_main_basesoc_rx_phase_cry_8_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(N_409_TMR_0),
    .S1(N_410_TMR_0)
  );
  defparam un5_main_basesoc_rx_phase_cry_7_0_TMR_0.INIT0 = "50AA";
  defparam un5_main_basesoc_rx_phase_cry_7_0_TMR_0.INIT1 = "50AA";
  defparam un5_main_basesoc_rx_phase_cry_7_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57141.8-57154.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_7_0_TMR_1 (
    .A0(dsp_join_kb_27_TMR_1[7]),
    .A1(dsp_join_kb_27_TMR_1[8]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(un5_main_basesoc_rx_phase_cry_6_TMR_1),
    .COUT(un5_main_basesoc_rx_phase_cry_8_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(N_409_TMR_1),
    .S1(N_410_TMR_1)
  );
  defparam un5_main_basesoc_rx_phase_cry_7_0_TMR_1.INIT0 = "50AA";
  defparam un5_main_basesoc_rx_phase_cry_7_0_TMR_1.INIT1 = "50AA";
  defparam un5_main_basesoc_rx_phase_cry_7_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57141.8-57154.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_7_0_TMR_2 (
    .A0(dsp_join_kb_27_TMR_2[7]),
    .A1(dsp_join_kb_27_TMR_2[8]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(un5_main_basesoc_rx_phase_cry_6_TMR_2),
    .COUT(un5_main_basesoc_rx_phase_cry_8_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(N_409_TMR_2),
    .S1(N_410_TMR_2)
  );
  defparam un5_main_basesoc_rx_phase_cry_7_0_TMR_2.INIT0 = "50AA";
  defparam un5_main_basesoc_rx_phase_cry_7_0_TMR_2.INIT1 = "50AA";
  defparam un5_main_basesoc_rx_phase_cry_7_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57123.8-57136.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_9_0_TMR_0 (
    .A0(dsp_join_kb_27_TMR_0[9]),
    .A1(dsp_join_kb_27_TMR_0[10]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(un5_main_basesoc_rx_phase_cry_8_TMR_0),
    .COUT(un5_main_basesoc_rx_phase_cry_10_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(N_411_TMR_0),
    .S1(N_412_TMR_0)
  );
  defparam un5_main_basesoc_rx_phase_cry_9_0_TMR_0.INIT0 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_9_0_TMR_0.INIT1 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_9_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57123.8-57136.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_9_0_TMR_1 (
    .A0(dsp_join_kb_27_TMR_1[9]),
    .A1(dsp_join_kb_27_TMR_1[10]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(un5_main_basesoc_rx_phase_cry_8_TMR_1),
    .COUT(un5_main_basesoc_rx_phase_cry_10_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(N_411_TMR_1),
    .S1(N_412_TMR_1)
  );
  defparam un5_main_basesoc_rx_phase_cry_9_0_TMR_1.INIT0 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_9_0_TMR_1.INIT1 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_9_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57123.8-57136.2" *)
  CCU2 un5_main_basesoc_rx_phase_cry_9_0_TMR_2 (
    .A0(dsp_join_kb_27_TMR_2[9]),
    .A1(dsp_join_kb_27_TMR_2[10]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(un5_main_basesoc_rx_phase_cry_8_TMR_2),
    .COUT(un5_main_basesoc_rx_phase_cry_10_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(N_411_TMR_2),
    .S1(N_412_TMR_2)
  );
  defparam un5_main_basesoc_rx_phase_cry_9_0_TMR_2.INIT0 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_9_0_TMR_2.INIT1 = "A033";
  defparam un5_main_basesoc_rx_phase_cry_9_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57517.8-57530.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_0_0_TMR_0 (
    .A0(VCC_TMR_0),
    .A1(dsp_join_kb_26_TMR_0[0]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(GND_0),
    .COUT(un5_main_basesoc_tx_phase_cry_0_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un5_main_basesoc_tx_phase_cry_0_0_S0_TMR_0),
    .S1(un5_main_basesoc_tx_phase_cry_0_0_S1_TMR_0)
  );
  defparam un5_main_basesoc_tx_phase_cry_0_0_TMR_0.INIT0 = "5033";
  defparam un5_main_basesoc_tx_phase_cry_0_0_TMR_0.INIT1 = "50AA";
  defparam un5_main_basesoc_tx_phase_cry_0_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57517.8-57530.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_0_0_TMR_1 (
    .A0(VCC_TMR_1),
    .A1(dsp_join_kb_26_TMR_1[0]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(GND_0),
    .COUT(un5_main_basesoc_tx_phase_cry_0_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un5_main_basesoc_tx_phase_cry_0_0_S0_TMR_1),
    .S1(un5_main_basesoc_tx_phase_cry_0_0_S1_TMR_1)
  );
  defparam un5_main_basesoc_tx_phase_cry_0_0_TMR_1.INIT0 = "5033";
  defparam un5_main_basesoc_tx_phase_cry_0_0_TMR_1.INIT1 = "50AA";
  defparam un5_main_basesoc_tx_phase_cry_0_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57517.8-57530.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_0_0_TMR_2 (
    .A0(VCC_TMR_2),
    .A1(dsp_join_kb_26_TMR_2[0]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(GND_0),
    .COUT(un5_main_basesoc_tx_phase_cry_0_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un5_main_basesoc_tx_phase_cry_0_0_S0_TMR_2),
    .S1(un5_main_basesoc_tx_phase_cry_0_0_S1_TMR_2)
  );
  defparam un5_main_basesoc_tx_phase_cry_0_0_TMR_2.INIT0 = "5033";
  defparam un5_main_basesoc_tx_phase_cry_0_0_TMR_2.INIT1 = "50AA";
  defparam un5_main_basesoc_tx_phase_cry_0_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57410.8-57423.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_11_0_TMR_0 (
    .A0(dsp_join_kb_26_TMR_0[11]),
    .A1(dsp_join_kb_26_TMR_0[12]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(un5_main_basesoc_tx_phase_cry_10_TMR_0),
    .COUT(un5_main_basesoc_tx_phase_cry_12_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un5_main_basesoc_tx_phase_cry_11_0_S0_TMR_0),
    .S1(un5_main_basesoc_tx_phase_cry_11_0_S1_TMR_0)
  );
  defparam un5_main_basesoc_tx_phase_cry_11_0_TMR_0.INIT0 = "50AA";
  defparam un5_main_basesoc_tx_phase_cry_11_0_TMR_0.INIT1 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_11_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57410.8-57423.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_11_0_TMR_1 (
    .A0(dsp_join_kb_26_TMR_1[11]),
    .A1(dsp_join_kb_26_TMR_1[12]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(un5_main_basesoc_tx_phase_cry_10_TMR_1),
    .COUT(un5_main_basesoc_tx_phase_cry_12_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un5_main_basesoc_tx_phase_cry_11_0_S0_TMR_1),
    .S1(un5_main_basesoc_tx_phase_cry_11_0_S1_TMR_1)
  );
  defparam un5_main_basesoc_tx_phase_cry_11_0_TMR_1.INIT0 = "50AA";
  defparam un5_main_basesoc_tx_phase_cry_11_0_TMR_1.INIT1 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_11_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57410.8-57423.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_11_0_TMR_2 (
    .A0(dsp_join_kb_26_TMR_2[11]),
    .A1(dsp_join_kb_26_TMR_2[12]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(un5_main_basesoc_tx_phase_cry_10_TMR_2),
    .COUT(un5_main_basesoc_tx_phase_cry_12_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un5_main_basesoc_tx_phase_cry_11_0_S0_TMR_2),
    .S1(un5_main_basesoc_tx_phase_cry_11_0_S1_TMR_2)
  );
  defparam un5_main_basesoc_tx_phase_cry_11_0_TMR_2.INIT0 = "50AA";
  defparam un5_main_basesoc_tx_phase_cry_11_0_TMR_2.INIT1 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_11_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57392.8-57405.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_13_0_TMR_0 (
    .A0(dsp_join_kb_26_TMR_0[13]),
    .A1(dsp_join_kb_26_TMR_0[14]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(un5_main_basesoc_tx_phase_cry_12_TMR_0),
    .COUT(un5_main_basesoc_tx_phase_cry_14_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un5_main_basesoc_tx_phase_cry_13_0_S0_TMR_0),
    .S1(un5_main_basesoc_tx_phase_cry_13_0_S1_TMR_0)
  );
  defparam un5_main_basesoc_tx_phase_cry_13_0_TMR_0.INIT0 = "50AA";
  defparam un5_main_basesoc_tx_phase_cry_13_0_TMR_0.INIT1 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_13_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57392.8-57405.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_13_0_TMR_1 (
    .A0(dsp_join_kb_26_TMR_1[13]),
    .A1(dsp_join_kb_26_TMR_1[14]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(un5_main_basesoc_tx_phase_cry_12_TMR_1),
    .COUT(un5_main_basesoc_tx_phase_cry_14_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un5_main_basesoc_tx_phase_cry_13_0_S0_TMR_1),
    .S1(un5_main_basesoc_tx_phase_cry_13_0_S1_TMR_1)
  );
  defparam un5_main_basesoc_tx_phase_cry_13_0_TMR_1.INIT0 = "50AA";
  defparam un5_main_basesoc_tx_phase_cry_13_0_TMR_1.INIT1 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_13_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57392.8-57405.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_13_0_TMR_2 (
    .A0(dsp_join_kb_26_TMR_2[13]),
    .A1(dsp_join_kb_26_TMR_2[14]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(un5_main_basesoc_tx_phase_cry_12_TMR_2),
    .COUT(un5_main_basesoc_tx_phase_cry_14_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un5_main_basesoc_tx_phase_cry_13_0_S0_TMR_2),
    .S1(un5_main_basesoc_tx_phase_cry_13_0_S1_TMR_2)
  );
  defparam un5_main_basesoc_tx_phase_cry_13_0_TMR_2.INIT0 = "50AA";
  defparam un5_main_basesoc_tx_phase_cry_13_0_TMR_2.INIT1 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_13_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57374.8-57387.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_15_0_TMR_0 (
    .A0(dsp_join_kb_26_TMR_0[15]),
    .A1(dsp_join_kb_26_TMR_0[16]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(un5_main_basesoc_tx_phase_cry_14_TMR_0),
    .COUT(un5_main_basesoc_tx_phase_cry_16_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un5_main_basesoc_tx_phase_cry_15_0_S0_TMR_0),
    .S1(un5_main_basesoc_tx_phase_cry_15_0_S1_TMR_0)
  );
  defparam un5_main_basesoc_tx_phase_cry_15_0_TMR_0.INIT0 = "50AA";
  defparam un5_main_basesoc_tx_phase_cry_15_0_TMR_0.INIT1 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_15_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57374.8-57387.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_15_0_TMR_1 (
    .A0(dsp_join_kb_26_TMR_1[15]),
    .A1(dsp_join_kb_26_TMR_1[16]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(un5_main_basesoc_tx_phase_cry_14_TMR_1),
    .COUT(un5_main_basesoc_tx_phase_cry_16_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un5_main_basesoc_tx_phase_cry_15_0_S0_TMR_1),
    .S1(un5_main_basesoc_tx_phase_cry_15_0_S1_TMR_1)
  );
  defparam un5_main_basesoc_tx_phase_cry_15_0_TMR_1.INIT0 = "50AA";
  defparam un5_main_basesoc_tx_phase_cry_15_0_TMR_1.INIT1 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_15_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57374.8-57387.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_15_0_TMR_2 (
    .A0(dsp_join_kb_26_TMR_2[15]),
    .A1(dsp_join_kb_26_TMR_2[16]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(un5_main_basesoc_tx_phase_cry_14_TMR_2),
    .COUT(un5_main_basesoc_tx_phase_cry_16_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un5_main_basesoc_tx_phase_cry_15_0_S0_TMR_2),
    .S1(un5_main_basesoc_tx_phase_cry_15_0_S1_TMR_2)
  );
  defparam un5_main_basesoc_tx_phase_cry_15_0_TMR_2.INIT0 = "50AA";
  defparam un5_main_basesoc_tx_phase_cry_15_0_TMR_2.INIT1 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_15_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57356.8-57369.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_17_0_TMR_0 (
    .A0(dsp_join_kb_26_TMR_0[17]),
    .A1(dsp_join_kb_26_TMR_0[18]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(un5_main_basesoc_tx_phase_cry_16_TMR_0),
    .COUT(un5_main_basesoc_tx_phase_cry_18_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un5_main_basesoc_tx_phase_cry_17_0_S0_TMR_0),
    .S1(un5_main_basesoc_tx_phase_cry_17_0_S1_TMR_0)
  );
  defparam un5_main_basesoc_tx_phase_cry_17_0_TMR_0.INIT0 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_17_0_TMR_0.INIT1 = "50AA";
  defparam un5_main_basesoc_tx_phase_cry_17_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57356.8-57369.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_17_0_TMR_1 (
    .A0(dsp_join_kb_26_TMR_1[17]),
    .A1(dsp_join_kb_26_TMR_1[18]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(un5_main_basesoc_tx_phase_cry_16_TMR_1),
    .COUT(un5_main_basesoc_tx_phase_cry_18_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un5_main_basesoc_tx_phase_cry_17_0_S0_TMR_1),
    .S1(un5_main_basesoc_tx_phase_cry_17_0_S1_TMR_1)
  );
  defparam un5_main_basesoc_tx_phase_cry_17_0_TMR_1.INIT0 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_17_0_TMR_1.INIT1 = "50AA";
  defparam un5_main_basesoc_tx_phase_cry_17_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57356.8-57369.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_17_0_TMR_2 (
    .A0(dsp_join_kb_26_TMR_2[17]),
    .A1(dsp_join_kb_26_TMR_2[18]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(un5_main_basesoc_tx_phase_cry_16_TMR_2),
    .COUT(un5_main_basesoc_tx_phase_cry_18_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un5_main_basesoc_tx_phase_cry_17_0_S0_TMR_2),
    .S1(un5_main_basesoc_tx_phase_cry_17_0_S1_TMR_2)
  );
  defparam un5_main_basesoc_tx_phase_cry_17_0_TMR_2.INIT0 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_17_0_TMR_2.INIT1 = "50AA";
  defparam un5_main_basesoc_tx_phase_cry_17_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57338.8-57351.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_19_0_TMR_0 (
    .A0(dsp_join_kb_26_TMR_0[19]),
    .A1(dsp_join_kb_26_TMR_0[20]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(un5_main_basesoc_tx_phase_cry_18_TMR_0),
    .COUT(un5_main_basesoc_tx_phase_cry_20_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un5_main_basesoc_tx_phase_cry_19_0_S0_TMR_0),
    .S1(un5_main_basesoc_tx_phase_cry_19_0_S1_TMR_0)
  );
  defparam un5_main_basesoc_tx_phase_cry_19_0_TMR_0.INIT0 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_19_0_TMR_0.INIT1 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_19_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57338.8-57351.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_19_0_TMR_1 (
    .A0(dsp_join_kb_26_TMR_1[19]),
    .A1(dsp_join_kb_26_TMR_1[20]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(un5_main_basesoc_tx_phase_cry_18_TMR_1),
    .COUT(un5_main_basesoc_tx_phase_cry_20_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un5_main_basesoc_tx_phase_cry_19_0_S0_TMR_1),
    .S1(un5_main_basesoc_tx_phase_cry_19_0_S1_TMR_1)
  );
  defparam un5_main_basesoc_tx_phase_cry_19_0_TMR_1.INIT0 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_19_0_TMR_1.INIT1 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_19_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57338.8-57351.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_19_0_TMR_2 (
    .A0(dsp_join_kb_26_TMR_2[19]),
    .A1(dsp_join_kb_26_TMR_2[20]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(un5_main_basesoc_tx_phase_cry_18_TMR_2),
    .COUT(un5_main_basesoc_tx_phase_cry_20_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un5_main_basesoc_tx_phase_cry_19_0_S0_TMR_2),
    .S1(un5_main_basesoc_tx_phase_cry_19_0_S1_TMR_2)
  );
  defparam un5_main_basesoc_tx_phase_cry_19_0_TMR_2.INIT0 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_19_0_TMR_2.INIT1 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_19_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57500.8-57513.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_1_0_TMR_0 (
    .A0(dsp_join_kb_26_TMR_0[1]),
    .A1(dsp_join_kb_26_TMR_0[2]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(un5_main_basesoc_tx_phase_cry_0_TMR_0),
    .COUT(un5_main_basesoc_tx_phase_cry_2_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un5_main_basesoc_tx_phase_cry_1_0_S0_TMR_0),
    .S1(un5_main_basesoc_tx_phase_cry_1_0_S1_TMR_0)
  );
  defparam un5_main_basesoc_tx_phase_cry_1_0_TMR_0.INIT0 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_1_0_TMR_0.INIT1 = "50AA";
  defparam un5_main_basesoc_tx_phase_cry_1_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57500.8-57513.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_1_0_TMR_1 (
    .A0(dsp_join_kb_26_TMR_1[1]),
    .A1(dsp_join_kb_26_TMR_1[2]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(un5_main_basesoc_tx_phase_cry_0_TMR_1),
    .COUT(un5_main_basesoc_tx_phase_cry_2_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un5_main_basesoc_tx_phase_cry_1_0_S0_TMR_1),
    .S1(un5_main_basesoc_tx_phase_cry_1_0_S1_TMR_1)
  );
  defparam un5_main_basesoc_tx_phase_cry_1_0_TMR_1.INIT0 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_1_0_TMR_1.INIT1 = "50AA";
  defparam un5_main_basesoc_tx_phase_cry_1_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57500.8-57513.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_1_0_TMR_2 (
    .A0(dsp_join_kb_26_TMR_2[1]),
    .A1(dsp_join_kb_26_TMR_2[2]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(un5_main_basesoc_tx_phase_cry_0_TMR_2),
    .COUT(un5_main_basesoc_tx_phase_cry_2_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un5_main_basesoc_tx_phase_cry_1_0_S0_TMR_2),
    .S1(un5_main_basesoc_tx_phase_cry_1_0_S1_TMR_2)
  );
  defparam un5_main_basesoc_tx_phase_cry_1_0_TMR_2.INIT0 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_1_0_TMR_2.INIT1 = "50AA";
  defparam un5_main_basesoc_tx_phase_cry_1_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57320.8-57333.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_21_0_TMR_0 (
    .A0(dsp_join_kb_26_TMR_0[21]),
    .A1(dsp_join_kb_26_TMR_0[22]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(un5_main_basesoc_tx_phase_cry_20_TMR_0),
    .COUT(un5_main_basesoc_tx_phase_cry_22_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un5_main_basesoc_tx_phase_cry_21_0_S0_TMR_0),
    .S1(un5_main_basesoc_tx_phase_cry_21_0_S1_TMR_0)
  );
  defparam un5_main_basesoc_tx_phase_cry_21_0_TMR_0.INIT0 = "50AA";
  defparam un5_main_basesoc_tx_phase_cry_21_0_TMR_0.INIT1 = "50AA";
  defparam un5_main_basesoc_tx_phase_cry_21_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57320.8-57333.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_21_0_TMR_1 (
    .A0(dsp_join_kb_26_TMR_1[21]),
    .A1(dsp_join_kb_26_TMR_1[22]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(un5_main_basesoc_tx_phase_cry_20_TMR_1),
    .COUT(un5_main_basesoc_tx_phase_cry_22_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un5_main_basesoc_tx_phase_cry_21_0_S0_TMR_1),
    .S1(un5_main_basesoc_tx_phase_cry_21_0_S1_TMR_1)
  );
  defparam un5_main_basesoc_tx_phase_cry_21_0_TMR_1.INIT0 = "50AA";
  defparam un5_main_basesoc_tx_phase_cry_21_0_TMR_1.INIT1 = "50AA";
  defparam un5_main_basesoc_tx_phase_cry_21_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57320.8-57333.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_21_0_TMR_2 (
    .A0(dsp_join_kb_26_TMR_2[21]),
    .A1(dsp_join_kb_26_TMR_2[22]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(un5_main_basesoc_tx_phase_cry_20_TMR_2),
    .COUT(un5_main_basesoc_tx_phase_cry_22_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un5_main_basesoc_tx_phase_cry_21_0_S0_TMR_2),
    .S1(un5_main_basesoc_tx_phase_cry_21_0_S1_TMR_2)
  );
  defparam un5_main_basesoc_tx_phase_cry_21_0_TMR_2.INIT0 = "50AA";
  defparam un5_main_basesoc_tx_phase_cry_21_0_TMR_2.INIT1 = "50AA";
  defparam un5_main_basesoc_tx_phase_cry_21_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57302.8-57315.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_23_0_TMR_0 (
    .A0(dsp_join_kb_26_TMR_0[23]),
    .A1(dsp_join_kb_26_TMR_0[24]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(un5_main_basesoc_tx_phase_cry_22_TMR_0),
    .COUT(un5_main_basesoc_tx_phase_cry_24_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un5_main_basesoc_tx_phase_cry_23_0_S0_TMR_0),
    .S1(un5_main_basesoc_tx_phase_cry_23_0_S1_TMR_0)
  );
  defparam un5_main_basesoc_tx_phase_cry_23_0_TMR_0.INIT0 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_23_0_TMR_0.INIT1 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_23_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57302.8-57315.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_23_0_TMR_1 (
    .A0(dsp_join_kb_26_TMR_1[23]),
    .A1(dsp_join_kb_26_TMR_1[24]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(un5_main_basesoc_tx_phase_cry_22_TMR_1),
    .COUT(un5_main_basesoc_tx_phase_cry_24_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un5_main_basesoc_tx_phase_cry_23_0_S0_TMR_1),
    .S1(un5_main_basesoc_tx_phase_cry_23_0_S1_TMR_1)
  );
  defparam un5_main_basesoc_tx_phase_cry_23_0_TMR_1.INIT0 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_23_0_TMR_1.INIT1 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_23_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57302.8-57315.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_23_0_TMR_2 (
    .A0(dsp_join_kb_26_TMR_2[23]),
    .A1(dsp_join_kb_26_TMR_2[24]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(un5_main_basesoc_tx_phase_cry_22_TMR_2),
    .COUT(un5_main_basesoc_tx_phase_cry_24_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un5_main_basesoc_tx_phase_cry_23_0_S0_TMR_2),
    .S1(un5_main_basesoc_tx_phase_cry_23_0_S1_TMR_2)
  );
  defparam un5_main_basesoc_tx_phase_cry_23_0_TMR_2.INIT0 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_23_0_TMR_2.INIT1 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_23_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57284.8-57297.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_25_0_TMR_0 (
    .A0(dsp_join_kb_26_TMR_0[25]),
    .A1(dsp_join_kb_26_TMR_0[26]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(un5_main_basesoc_tx_phase_cry_24_TMR_0),
    .COUT(un5_main_basesoc_tx_phase_cry_26_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un5_main_basesoc_tx_phase_cry_25_0_S0_TMR_0),
    .S1(un5_main_basesoc_tx_phase_cry_25_0_S1_TMR_0)
  );
  defparam un5_main_basesoc_tx_phase_cry_25_0_TMR_0.INIT0 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_25_0_TMR_0.INIT1 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_25_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57284.8-57297.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_25_0_TMR_1 (
    .A0(dsp_join_kb_26_TMR_1[25]),
    .A1(dsp_join_kb_26_TMR_1[26]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(un5_main_basesoc_tx_phase_cry_24_TMR_1),
    .COUT(un5_main_basesoc_tx_phase_cry_26_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un5_main_basesoc_tx_phase_cry_25_0_S0_TMR_1),
    .S1(un5_main_basesoc_tx_phase_cry_25_0_S1_TMR_1)
  );
  defparam un5_main_basesoc_tx_phase_cry_25_0_TMR_1.INIT0 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_25_0_TMR_1.INIT1 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_25_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57284.8-57297.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_25_0_TMR_2 (
    .A0(dsp_join_kb_26_TMR_2[25]),
    .A1(dsp_join_kb_26_TMR_2[26]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(un5_main_basesoc_tx_phase_cry_24_TMR_2),
    .COUT(un5_main_basesoc_tx_phase_cry_26_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un5_main_basesoc_tx_phase_cry_25_0_S0_TMR_2),
    .S1(un5_main_basesoc_tx_phase_cry_25_0_S1_TMR_2)
  );
  defparam un5_main_basesoc_tx_phase_cry_25_0_TMR_2.INIT0 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_25_0_TMR_2.INIT1 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_25_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57266.8-57279.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_27_0_TMR_0 (
    .A0(dsp_join_kb_26_TMR_0[27]),
    .A1(dsp_join_kb_26_TMR_0[28]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(un5_main_basesoc_tx_phase_cry_26_TMR_0),
    .COUT(un5_main_basesoc_tx_phase_cry_28_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un5_main_basesoc_tx_phase_cry_27_0_S0_TMR_0),
    .S1(un5_main_basesoc_tx_phase_cry_27_0_S1_TMR_0)
  );
  defparam un5_main_basesoc_tx_phase_cry_27_0_TMR_0.INIT0 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_27_0_TMR_0.INIT1 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_27_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57266.8-57279.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_27_0_TMR_1 (
    .A0(dsp_join_kb_26_TMR_1[27]),
    .A1(dsp_join_kb_26_TMR_1[28]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(un5_main_basesoc_tx_phase_cry_26_TMR_1),
    .COUT(un5_main_basesoc_tx_phase_cry_28_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un5_main_basesoc_tx_phase_cry_27_0_S0_TMR_1),
    .S1(un5_main_basesoc_tx_phase_cry_27_0_S1_TMR_1)
  );
  defparam un5_main_basesoc_tx_phase_cry_27_0_TMR_1.INIT0 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_27_0_TMR_1.INIT1 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_27_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57266.8-57279.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_27_0_TMR_2 (
    .A0(dsp_join_kb_26_TMR_2[27]),
    .A1(dsp_join_kb_26_TMR_2[28]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(un5_main_basesoc_tx_phase_cry_26_TMR_2),
    .COUT(un5_main_basesoc_tx_phase_cry_28_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un5_main_basesoc_tx_phase_cry_27_0_S0_TMR_2),
    .S1(un5_main_basesoc_tx_phase_cry_27_0_S1_TMR_2)
  );
  defparam un5_main_basesoc_tx_phase_cry_27_0_TMR_2.INIT0 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_27_0_TMR_2.INIT1 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_27_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57248.8-57261.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_29_0_TMR_0 (
    .A0(dsp_join_kb_26_TMR_0[29]),
    .A1(dsp_join_kb_26_TMR_0[30]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(un5_main_basesoc_tx_phase_cry_28_TMR_0),
    .COUT(un5_main_basesoc_tx_phase_cry_30_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un5_main_basesoc_tx_phase_cry_29_0_S0_TMR_0),
    .S1(un5_main_basesoc_tx_phase_cry_29_0_S1_TMR_0)
  );
  defparam un5_main_basesoc_tx_phase_cry_29_0_TMR_0.INIT0 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_29_0_TMR_0.INIT1 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_29_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57248.8-57261.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_29_0_TMR_1 (
    .A0(dsp_join_kb_26_TMR_1[29]),
    .A1(dsp_join_kb_26_TMR_1[30]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(un5_main_basesoc_tx_phase_cry_28_TMR_1),
    .COUT(un5_main_basesoc_tx_phase_cry_30_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un5_main_basesoc_tx_phase_cry_29_0_S0_TMR_1),
    .S1(un5_main_basesoc_tx_phase_cry_29_0_S1_TMR_1)
  );
  defparam un5_main_basesoc_tx_phase_cry_29_0_TMR_1.INIT0 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_29_0_TMR_1.INIT1 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_29_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57248.8-57261.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_29_0_TMR_2 (
    .A0(dsp_join_kb_26_TMR_2[29]),
    .A1(dsp_join_kb_26_TMR_2[30]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(un5_main_basesoc_tx_phase_cry_28_TMR_2),
    .COUT(un5_main_basesoc_tx_phase_cry_30_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un5_main_basesoc_tx_phase_cry_29_0_S0_TMR_2),
    .S1(un5_main_basesoc_tx_phase_cry_29_0_S1_TMR_2)
  );
  defparam un5_main_basesoc_tx_phase_cry_29_0_TMR_2.INIT0 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_29_0_TMR_2.INIT1 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_29_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57230.8-57243.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_31_0_TMR_0 (
    .A0(dsp_join_kb_26_TMR_0[31]),
    .A1(VCC_TMR_0),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(un5_main_basesoc_tx_phase_cry_30_TMR_0),
    .COUT(un5_main_basesoc_tx_phase_cry_31_0_COUT_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un5_main_basesoc_tx_phase_cry_31_0_S0_TMR_0),
    .S1(un5_main_basesoc_tx_phase_cry_31_TMR_0)
  );
  defparam un5_main_basesoc_tx_phase_cry_31_0_TMR_0.INIT0 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_31_0_TMR_0.INIT1 = "5033";
  defparam un5_main_basesoc_tx_phase_cry_31_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57230.8-57243.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_31_0_TMR_1 (
    .A0(dsp_join_kb_26_TMR_1[31]),
    .A1(VCC_TMR_1),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(un5_main_basesoc_tx_phase_cry_30_TMR_1),
    .COUT(un5_main_basesoc_tx_phase_cry_31_0_COUT_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un5_main_basesoc_tx_phase_cry_31_0_S0_TMR_1),
    .S1(un5_main_basesoc_tx_phase_cry_31_TMR_1)
  );
  defparam un5_main_basesoc_tx_phase_cry_31_0_TMR_1.INIT0 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_31_0_TMR_1.INIT1 = "5033";
  defparam un5_main_basesoc_tx_phase_cry_31_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57230.8-57243.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_31_0_TMR_2 (
    .A0(dsp_join_kb_26_TMR_2[31]),
    .A1(VCC_TMR_2),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(un5_main_basesoc_tx_phase_cry_30_TMR_2),
    .COUT(un5_main_basesoc_tx_phase_cry_31_0_COUT_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un5_main_basesoc_tx_phase_cry_31_0_S0_TMR_2),
    .S1(un5_main_basesoc_tx_phase_cry_31_TMR_2)
  );
  defparam un5_main_basesoc_tx_phase_cry_31_0_TMR_2.INIT0 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_31_0_TMR_2.INIT1 = "5033";
  defparam un5_main_basesoc_tx_phase_cry_31_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57482.8-57495.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_3_0_TMR_0 (
    .A0(dsp_join_kb_26_TMR_0[3]),
    .A1(dsp_join_kb_26_TMR_0[4]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(un5_main_basesoc_tx_phase_cry_2_TMR_0),
    .COUT(un5_main_basesoc_tx_phase_cry_4_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un5_main_basesoc_tx_phase_cry_3_0_S0_TMR_0),
    .S1(un5_main_basesoc_tx_phase_cry_3_0_S1_TMR_0)
  );
  defparam un5_main_basesoc_tx_phase_cry_3_0_TMR_0.INIT0 = "50AA";
  defparam un5_main_basesoc_tx_phase_cry_3_0_TMR_0.INIT1 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_3_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57482.8-57495.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_3_0_TMR_1 (
    .A0(dsp_join_kb_26_TMR_1[3]),
    .A1(dsp_join_kb_26_TMR_1[4]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(un5_main_basesoc_tx_phase_cry_2_TMR_1),
    .COUT(un5_main_basesoc_tx_phase_cry_4_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un5_main_basesoc_tx_phase_cry_3_0_S0_TMR_1),
    .S1(un5_main_basesoc_tx_phase_cry_3_0_S1_TMR_1)
  );
  defparam un5_main_basesoc_tx_phase_cry_3_0_TMR_1.INIT0 = "50AA";
  defparam un5_main_basesoc_tx_phase_cry_3_0_TMR_1.INIT1 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_3_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57482.8-57495.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_3_0_TMR_2 (
    .A0(dsp_join_kb_26_TMR_2[3]),
    .A1(dsp_join_kb_26_TMR_2[4]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(un5_main_basesoc_tx_phase_cry_2_TMR_2),
    .COUT(un5_main_basesoc_tx_phase_cry_4_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un5_main_basesoc_tx_phase_cry_3_0_S0_TMR_2),
    .S1(un5_main_basesoc_tx_phase_cry_3_0_S1_TMR_2)
  );
  defparam un5_main_basesoc_tx_phase_cry_3_0_TMR_2.INIT0 = "50AA";
  defparam un5_main_basesoc_tx_phase_cry_3_0_TMR_2.INIT1 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_3_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57464.8-57477.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_5_0_TMR_0 (
    .A0(dsp_join_kb_26_TMR_0[5]),
    .A1(dsp_join_kb_26_TMR_0[6]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(un5_main_basesoc_tx_phase_cry_4_TMR_0),
    .COUT(un5_main_basesoc_tx_phase_cry_6_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un5_main_basesoc_tx_phase_cry_5_0_S0_TMR_0),
    .S1(un5_main_basesoc_tx_phase_cry_5_0_S1_TMR_0)
  );
  defparam un5_main_basesoc_tx_phase_cry_5_0_TMR_0.INIT0 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_5_0_TMR_0.INIT1 = "50AA";
  defparam un5_main_basesoc_tx_phase_cry_5_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57464.8-57477.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_5_0_TMR_1 (
    .A0(dsp_join_kb_26_TMR_1[5]),
    .A1(dsp_join_kb_26_TMR_1[6]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(un5_main_basesoc_tx_phase_cry_4_TMR_1),
    .COUT(un5_main_basesoc_tx_phase_cry_6_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un5_main_basesoc_tx_phase_cry_5_0_S0_TMR_1),
    .S1(un5_main_basesoc_tx_phase_cry_5_0_S1_TMR_1)
  );
  defparam un5_main_basesoc_tx_phase_cry_5_0_TMR_1.INIT0 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_5_0_TMR_1.INIT1 = "50AA";
  defparam un5_main_basesoc_tx_phase_cry_5_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57464.8-57477.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_5_0_TMR_2 (
    .A0(dsp_join_kb_26_TMR_2[5]),
    .A1(dsp_join_kb_26_TMR_2[6]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(un5_main_basesoc_tx_phase_cry_4_TMR_2),
    .COUT(un5_main_basesoc_tx_phase_cry_6_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un5_main_basesoc_tx_phase_cry_5_0_S0_TMR_2),
    .S1(un5_main_basesoc_tx_phase_cry_5_0_S1_TMR_2)
  );
  defparam un5_main_basesoc_tx_phase_cry_5_0_TMR_2.INIT0 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_5_0_TMR_2.INIT1 = "50AA";
  defparam un5_main_basesoc_tx_phase_cry_5_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57446.8-57459.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_7_0_TMR_0 (
    .A0(dsp_join_kb_26_TMR_0[7]),
    .A1(dsp_join_kb_26_TMR_0[8]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(un5_main_basesoc_tx_phase_cry_6_TMR_0),
    .COUT(un5_main_basesoc_tx_phase_cry_8_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un5_main_basesoc_tx_phase_cry_7_0_S0_TMR_0),
    .S1(un5_main_basesoc_tx_phase_cry_7_0_S1_TMR_0)
  );
  defparam un5_main_basesoc_tx_phase_cry_7_0_TMR_0.INIT0 = "50AA";
  defparam un5_main_basesoc_tx_phase_cry_7_0_TMR_0.INIT1 = "50AA";
  defparam un5_main_basesoc_tx_phase_cry_7_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57446.8-57459.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_7_0_TMR_1 (
    .A0(dsp_join_kb_26_TMR_1[7]),
    .A1(dsp_join_kb_26_TMR_1[8]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(un5_main_basesoc_tx_phase_cry_6_TMR_1),
    .COUT(un5_main_basesoc_tx_phase_cry_8_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un5_main_basesoc_tx_phase_cry_7_0_S0_TMR_1),
    .S1(un5_main_basesoc_tx_phase_cry_7_0_S1_TMR_1)
  );
  defparam un5_main_basesoc_tx_phase_cry_7_0_TMR_1.INIT0 = "50AA";
  defparam un5_main_basesoc_tx_phase_cry_7_0_TMR_1.INIT1 = "50AA";
  defparam un5_main_basesoc_tx_phase_cry_7_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57446.8-57459.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_7_0_TMR_2 (
    .A0(dsp_join_kb_26_TMR_2[7]),
    .A1(dsp_join_kb_26_TMR_2[8]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(un5_main_basesoc_tx_phase_cry_6_TMR_2),
    .COUT(un5_main_basesoc_tx_phase_cry_8_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un5_main_basesoc_tx_phase_cry_7_0_S0_TMR_2),
    .S1(un5_main_basesoc_tx_phase_cry_7_0_S1_TMR_2)
  );
  defparam un5_main_basesoc_tx_phase_cry_7_0_TMR_2.INIT0 = "50AA";
  defparam un5_main_basesoc_tx_phase_cry_7_0_TMR_2.INIT1 = "50AA";
  defparam un5_main_basesoc_tx_phase_cry_7_0_TMR_2.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57428.8-57441.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_9_0_TMR_0 (
    .A0(dsp_join_kb_26_TMR_0[9]),
    .A1(dsp_join_kb_26_TMR_0[10]),
    .B0(VCC_TMR_0),
    .B1(VCC_TMR_0),
    .C0(VCC_TMR_0),
    .C1(VCC_TMR_0),
    .CIN(un5_main_basesoc_tx_phase_cry_8_TMR_0),
    .COUT(un5_main_basesoc_tx_phase_cry_10_TMR_0),
    .D0(VCC_TMR_0),
    .D1(VCC_TMR_0),
    .S0(un5_main_basesoc_tx_phase_cry_9_0_S0_TMR_0),
    .S1(un5_main_basesoc_tx_phase_cry_9_0_S1_TMR_0)
  );
  defparam un5_main_basesoc_tx_phase_cry_9_0_TMR_0.INIT0 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_9_0_TMR_0.INIT1 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_9_0_TMR_0.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57428.8-57441.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_9_0_TMR_1 (
    .A0(dsp_join_kb_26_TMR_1[9]),
    .A1(dsp_join_kb_26_TMR_1[10]),
    .B0(VCC_TMR_1),
    .B1(VCC_TMR_1),
    .C0(VCC_TMR_1),
    .C1(VCC_TMR_1),
    .CIN(un5_main_basesoc_tx_phase_cry_8_TMR_1),
    .COUT(un5_main_basesoc_tx_phase_cry_10_TMR_1),
    .D0(VCC_TMR_1),
    .D1(VCC_TMR_1),
    .S0(un5_main_basesoc_tx_phase_cry_9_0_S0_TMR_1),
    .S1(un5_main_basesoc_tx_phase_cry_9_0_S1_TMR_1)
  );
  defparam un5_main_basesoc_tx_phase_cry_9_0_TMR_1.INIT0 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_9_0_TMR_1.INIT1 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_9_0_TMR_1.INJECT = "NO";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:57428.8-57441.2" *)
  CCU2 un5_main_basesoc_tx_phase_cry_9_0_TMR_2 (
    .A0(dsp_join_kb_26_TMR_2[9]),
    .A1(dsp_join_kb_26_TMR_2[10]),
    .B0(VCC_TMR_2),
    .B1(VCC_TMR_2),
    .C0(VCC_TMR_2),
    .C1(VCC_TMR_2),
    .CIN(un5_main_basesoc_tx_phase_cry_8_TMR_2),
    .COUT(un5_main_basesoc_tx_phase_cry_10_TMR_2),
    .D0(VCC_TMR_2),
    .D1(VCC_TMR_2),
    .S0(un5_main_basesoc_tx_phase_cry_9_0_S0_TMR_2),
    .S1(un5_main_basesoc_tx_phase_cry_9_0_S1_TMR_2)
  );
  defparam un5_main_basesoc_tx_phase_cry_9_0_TMR_2.INIT0 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_9_0_TMR_2.INIT1 = "A033";
  defparam un5_main_basesoc_tx_phase_cry_9_0_TMR_2.INJECT = "NO";
  LUT4 user_led0_c_0_RED_VOTER (
    .A(user_led0_c_TMR_0),
    .B(user_led0_c_TMR_1),
    .C(user_led0_c_TMR_2),
    .D(1'h0),
    .Z(user_led0_c_0_RED_VOTER_wire)
  );
  defparam user_led0_c_0_RED_VOTER.INIT = "0xFCC0";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55558.6-55561.2" *)
  OB user_led0_pad (
    .I(user_led0_c_0_RED_VOTER_wire),
    .O(user_led0)
  );
  LUT4 user_led10_c_0_RED_VOTER (
    .A(user_led10_c_TMR_0),
    .B(user_led10_c_TMR_1),
    .C(user_led10_c_TMR_2),
    .D(1'h0),
    .Z(user_led10_c_0_RED_VOTER_wire)
  );
  defparam user_led10_c_0_RED_VOTER.INIT = "0xFCC0";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55508.6-55511.2" *)
  OB user_led10_pad (
    .I(user_led10_c_0_RED_VOTER_wire),
    .O(user_led10)
  );
  LUT4 user_led11_c_0_RED_VOTER (
    .A(user_led11_c_TMR_0),
    .B(user_led11_c_TMR_1),
    .C(user_led11_c_TMR_2),
    .D(1'h0),
    .Z(user_led11_c_0_RED_VOTER_wire)
  );
  defparam user_led11_c_0_RED_VOTER.INIT = "0xFCC0";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55503.6-55506.2" *)
  OB user_led11_pad (
    .I(user_led11_c_0_RED_VOTER_wire),
    .O(user_led11)
  );
  LUT4 user_led12_c_0_RED_VOTER (
    .A(user_led12_c_TMR_0),
    .B(user_led12_c_TMR_1),
    .C(user_led12_c_TMR_2),
    .D(1'h0),
    .Z(user_led12_c_0_RED_VOTER_wire)
  );
  defparam user_led12_c_0_RED_VOTER.INIT = "0xFCC0";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55498.6-55501.2" *)
  OB user_led12_pad (
    .I(user_led12_c_0_RED_VOTER_wire),
    .O(user_led12)
  );
  LUT4 user_led13_c_0_RED_VOTER (
    .A(user_led13_c_TMR_0),
    .B(user_led13_c_TMR_1),
    .C(user_led13_c_TMR_2),
    .D(1'h0),
    .Z(user_led13_c_0_RED_VOTER_wire)
  );
  defparam user_led13_c_0_RED_VOTER.INIT = "0xFCC0";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55493.6-55496.2" *)
  OB user_led13_pad (
    .I(user_led13_c_0_RED_VOTER_wire),
    .O(user_led13)
  );
  LUT4 user_led1_c_0_RED_VOTER (
    .A(user_led1_c_TMR_0),
    .B(user_led1_c_TMR_1),
    .C(user_led1_c_TMR_2),
    .D(1'h0),
    .Z(user_led1_c_0_RED_VOTER_wire)
  );
  defparam user_led1_c_0_RED_VOTER.INIT = "0xFCC0";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55553.6-55556.2" *)
  OB user_led1_pad (
    .I(user_led1_c_0_RED_VOTER_wire),
    .O(user_led1)
  );
  LUT4 user_led2_c_0_RED_VOTER (
    .A(user_led2_c_TMR_0),
    .B(user_led2_c_TMR_1),
    .C(user_led2_c_TMR_2),
    .D(1'h0),
    .Z(user_led2_c_0_RED_VOTER_wire)
  );
  defparam user_led2_c_0_RED_VOTER.INIT = "0xFCC0";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55548.6-55551.2" *)
  OB user_led2_pad (
    .I(user_led2_c_0_RED_VOTER_wire),
    .O(user_led2)
  );
  LUT4 user_led3_c_0_RED_VOTER (
    .A(user_led3_c_TMR_0),
    .B(user_led3_c_TMR_1),
    .C(user_led3_c_TMR_2),
    .D(1'h0),
    .Z(user_led3_c_0_RED_VOTER_wire)
  );
  defparam user_led3_c_0_RED_VOTER.INIT = "0xFCC0";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55543.6-55546.2" *)
  OB user_led3_pad (
    .I(user_led3_c_0_RED_VOTER_wire),
    .O(user_led3)
  );
  LUT4 user_led4_c_0_RED_VOTER (
    .A(user_led4_c_TMR_0),
    .B(user_led4_c_TMR_1),
    .C(user_led4_c_TMR_2),
    .D(1'h0),
    .Z(user_led4_c_0_RED_VOTER_wire)
  );
  defparam user_led4_c_0_RED_VOTER.INIT = "0xFCC0";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55538.6-55541.2" *)
  OB user_led4_pad (
    .I(user_led4_c_0_RED_VOTER_wire),
    .O(user_led4)
  );
  LUT4 user_led5_c_0_RED_VOTER (
    .A(user_led5_c_TMR_0),
    .B(user_led5_c_TMR_1),
    .C(user_led5_c_TMR_2),
    .D(1'h0),
    .Z(user_led5_c_0_RED_VOTER_wire)
  );
  defparam user_led5_c_0_RED_VOTER.INIT = "0xFCC0";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55533.6-55536.2" *)
  OB user_led5_pad (
    .I(user_led5_c_0_RED_VOTER_wire),
    .O(user_led5)
  );
  LUT4 user_led6_c_0_RED_VOTER (
    .A(user_led6_c_TMR_0),
    .B(user_led6_c_TMR_1),
    .C(user_led6_c_TMR_2),
    .D(1'h0),
    .Z(user_led6_c_0_RED_VOTER_wire)
  );
  defparam user_led6_c_0_RED_VOTER.INIT = "0xFCC0";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55528.6-55531.2" *)
  OB user_led6_pad (
    .I(user_led6_c_0_RED_VOTER_wire),
    .O(user_led6)
  );
  LUT4 user_led7_c_0_RED_VOTER (
    .A(user_led7_c_TMR_0),
    .B(user_led7_c_TMR_1),
    .C(user_led7_c_TMR_2),
    .D(1'h0),
    .Z(user_led7_c_0_RED_VOTER_wire)
  );
  defparam user_led7_c_0_RED_VOTER.INIT = "0xFCC0";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55523.6-55526.2" *)
  OB user_led7_pad (
    .I(user_led7_c_0_RED_VOTER_wire),
    .O(user_led7)
  );
  LUT4 user_led8_c_0_RED_VOTER (
    .A(user_led8_c_TMR_0),
    .B(user_led8_c_TMR_1),
    .C(user_led8_c_TMR_2),
    .D(1'h0),
    .Z(user_led8_c_0_RED_VOTER_wire)
  );
  defparam user_led8_c_0_RED_VOTER.INIT = "0xFCC0";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55518.6-55521.2" *)
  OB user_led8_pad (
    .I(user_led8_c_0_RED_VOTER_wire),
    .O(user_led8)
  );
  LUT4 user_led9_c_0_RED_VOTER (
    .A(user_led9_c_TMR_0),
    .B(user_led9_c_TMR_1),
    .C(user_led9_c_TMR_2),
    .D(1'h0),
    .Z(user_led9_c_0_RED_VOTER_wire)
  );
  defparam user_led9_c_0_RED_VOTER.INIT = "0xFCC0";
  (* module_not_derived = 32'd1 *)
  (* src = "lattice_riscv.v:55513.6-55516.2" *)
  OB user_led9_pad (
    .I(user_led9_c_0_RED_VOTER_wire),
    .O(user_led9)
  );
endmodule
