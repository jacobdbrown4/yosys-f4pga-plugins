//Generated from netlist by SpyDrNet
//netlist name: zpu_core
module zpu_core
(
    areset,
    break,
    clk,
    enable,
    in_mem_busy,
    interrupt,
    out_mem_readEnable,
    out_mem_writeEnable,
    .mem_read[31:0]({mem_read[31], mem_read[30], mem_read[29], mem_read[28], mem_read[27], mem_read[26], mem_read[25], mem_read[24], mem_read[23], mem_read[22], mem_read[21], mem_read[20], mem_read[19], mem_read[18], mem_read[17], mem_read[16], mem_read[15], mem_read[14], mem_read[13], mem_read[12], mem_read[11], mem_read[10], mem_read[9], mem_read[8], mem_read[7], mem_read[6], mem_read[5], mem_read[4], mem_read[3], mem_read[2], mem_read[1], mem_read[0]}),
    .mem_write[31:0]({mem_write[31], mem_write[30], mem_write[29], mem_write[28], mem_write[27], mem_write[26], mem_write[25], mem_write[24], mem_write[23], mem_write[22], mem_write[21], mem_write[20], mem_write[19], mem_write[18], mem_write[17], mem_write[16], mem_write[15], mem_write[14], mem_write[13], mem_write[12], mem_write[11], mem_write[10], mem_write[9], mem_write[8], mem_write[7], mem_write[6], mem_write[5], mem_write[4], mem_write[3], mem_write[2], mem_write[1], mem_write[0]}),
    .mem_writeMask[3:0]({mem_writeMask[3], mem_writeMask[2], mem_writeMask[1], mem_writeMask[0]}),
    .out_mem_addr[15:0]({out_mem_addr[15], out_mem_addr[14], out_mem_addr[13], out_mem_addr[12], out_mem_addr[11], out_mem_addr[10], out_mem_addr[9], out_mem_addr[8], out_mem_addr[7], out_mem_addr[6], out_mem_addr[5], out_mem_addr[4], out_mem_addr[3], out_mem_addr[2], out_mem_addr[1], out_mem_addr[0]})
);

    input areset;
    output break;
    input clk;
    input enable;
    input in_mem_busy;
    input interrupt;
    output out_mem_readEnable;
    output out_mem_writeEnable;
    input [31:0]mem_read;
    output [31:0]mem_write;
    output [3:0]mem_writeMask;
    output [15:0]out_mem_addr;

    wire <const0>;
    wire <const1>;
    wire FSM_sequential_state[0]_i_1_n_0;
    wire FSM_sequential_state[0]_i_2_n_0;
    wire FSM_sequential_state[0]_i_3_n_0;
    wire FSM_sequential_state[0]_i_4_n_0;
    wire FSM_sequential_state[0]_i_5_n_0;
    wire FSM_sequential_state[0]_i_6_n_0;
    wire FSM_sequential_state[1]_i_3_n_0;
    wire FSM_sequential_state[2]_i_3_n_0;
    wire FSM_sequential_state[3]_i_1_n_0;
    wire FSM_sequential_state[3]_i_3_n_0;
    wire FSM_sequential_state[3]_i_5_n_0;
    wire [3:0]FSM_sequential_state_reg_n_0_;
    wire areset;
    wire areset_IBUF;
    wire break;
    wire break_OBUF;
    wire break_i_1_n_0;
    wire break_i_2_n_0;
    wire clk;
    wire clk_IBUF;
    wire clk_IBUF_BUFG;
    wire [1:0]data0;
    wire [14:1]data2;
    wire [4:0]decodedOpcode;
    wire decodedOpcode[4]_i_2_n_0;
    wire decodedOpcode[4]_i_5_n_0;
    wire [4:0]decodedOpcode_reg_n_0_;
    wire g0_b0__0_n_0;
    wire g0_b0_n_0;
    wire idim_flag;
    wire idim_flag_i_1_n_0;
    wire inInterrupt_i_1_n_0;
    wire inInterrupt_reg_n_0;
    wire in_mem_busy;
    wire in_mem_busy_IBUF;
    wire interrupt;
    wire interrupt_IBUF;
    wire [14:2]memAAddr;
    wire memAAddr[10]_i_4_n_0;
    wire memAAddr[11]_i_4_n_0;
    wire memAAddr[12]_i_4_n_0;
    wire memAAddr[13]_i_4_n_0;
    wire memAAddr[14]_i_4_n_0;
    wire memAAddr[14]_i_5_n_0;
    wire memAAddr[14]_i_6_n_0;
    wire memAAddr[2]_i_3_n_0;
    wire memAAddr[2]_i_4_n_0;
    wire memAAddr[3]_i_4_n_0;
    wire memAAddr[4]_i_4_n_0;
    wire memAAddr[5]_i_4_n_0;
    wire memAAddr[6]_i_4_n_0;
    wire memAAddr[7]_i_4_n_0;
    wire memAAddr[8]_i_4_n_0;
    wire memAAddr[9]_i_4_n_0;
    wire [14:2]memAAddr_reg_n_0_;
    wire [31:0]memARead;
    wire memAWriteEnable;
    wire memAWriteEnable_reg_n_0;
    wire [31:0]memAWrite;
    wire memAWrite[0]_i_4_n_0;
    wire memAWrite[10]_i_4_n_0;
    wire memAWrite[10]_i_7_n_0;
    wire memAWrite[11]_i_4_n_0;
    wire memAWrite[11]_i_7_n_0;
    wire memAWrite[12]_i_4_n_0;
    wire memAWrite[12]_i_7_n_0;
    wire memAWrite[13]_i_4_n_0;
    wire memAWrite[13]_i_7_n_0;
    wire memAWrite[14]_i_4_n_0;
    wire memAWrite[14]_i_7_n_0;
    wire memAWrite[1]_i_4_n_0;
    wire memAWrite[2]_i_4_n_0;
    wire memAWrite[2]_i_5_n_0;
    wire memAWrite[31]_i_4_n_0;
    wire memAWrite[3]_i_4_n_0;
    wire memAWrite[3]_i_5_n_0;
    wire memAWrite[4]_i_4_n_0;
    wire memAWrite[4]_i_5_n_0;
    wire memAWrite[5]_i_4_n_0;
    wire memAWrite[5]_i_5_n_0;
    wire memAWrite[6]_i_4_n_0;
    wire memAWrite[6]_i_5_n_0;
    wire memAWrite[7]_i_4_n_0;
    wire memAWrite[7]_i_7_n_0;
    wire memAWrite[8]_i_4_n_0;
    wire memAWrite[8]_i_7_n_0;
    wire memAWrite[9]_i_4_n_0;
    wire memAWrite[9]_i_7_n_0;
    wire [31:0]memAWrite_reg_n_0_;
    wire [14:2]memBAddr;
    wire memBAddr[13]_i_3_n_0;
    wire memBAddr[13]_i_4_n_0;
    wire memBAddr[13]_i_5_n_0;
    wire memBAddr[13]_i_6_n_0;
    wire memBAddr[14]_i_3_n_0;
    wire memBAddr[5]_i_3_n_0;
    wire memBAddr[5]_i_4_n_0;
    wire memBAddr[5]_i_5_n_0;
    wire memBAddr[5]_i_6_n_0;
    wire memBAddr[9]_i_3_n_0;
    wire memBAddr[9]_i_4_n_0;
    wire memBAddr[9]_i_5_n_0;
    wire memBAddr[9]_i_6_n_0;
    wire memBAddr_reg[13]_i_2_n_0;
    wire memBAddr_reg[13]_i_2_n_1;
    wire memBAddr_reg[13]_i_2_n_2;
    wire memBAddr_reg[13]_i_2_n_3;
    wire memBAddr_reg[13]_i_2_n_4;
    wire memBAddr_reg[13]_i_2_n_5;
    wire memBAddr_reg[13]_i_2_n_6;
    wire memBAddr_reg[13]_i_2_n_7;
    wire memBAddr_reg[14]_i_2_n_7;
    wire memBAddr_reg[5]_i_2_n_0;
    wire memBAddr_reg[5]_i_2_n_1;
    wire memBAddr_reg[5]_i_2_n_2;
    wire memBAddr_reg[5]_i_2_n_3;
    wire memBAddr_reg[5]_i_2_n_4;
    wire memBAddr_reg[5]_i_2_n_5;
    wire memBAddr_reg[5]_i_2_n_6;
    wire memBAddr_reg[5]_i_2_n_7;
    wire memBAddr_reg[9]_i_2_n_0;
    wire memBAddr_reg[9]_i_2_n_1;
    wire memBAddr_reg[9]_i_2_n_2;
    wire memBAddr_reg[9]_i_2_n_3;
    wire memBAddr_reg[9]_i_2_n_4;
    wire memBAddr_reg[9]_i_2_n_5;
    wire memBAddr_reg[9]_i_2_n_6;
    wire memBAddr_reg[9]_i_2_n_7;
    wire [14:2]memBAddr_reg_n_0_;
    wire [31:0]memBRead;
    wire memBWriteEnable;
    wire memBWriteEnable_reg_n_0;
    wire [31:0]memBWrite;
    wire [31:0]mem_read;
    wire [31:0]mem_read_IBUF;
    wire [3:0]mem_writeMask;
    wire [31:0]mem_write;
    wire mem_write[31]_i_1_n_0;
    wire [31:0]mem_write_OBUF;
    wire memory_n_0;
    wire memory_n_1;
    wire memory_n_148;
    wire memory_n_149;
    wire memory_n_150;
    wire memory_n_151;
    wire memory_n_152;
    wire memory_n_2;
    wire memory_n_3;
    wire memory_n_41;
    wire memory_n_42;
    wire [6:0]opcode_reg_n_0_;
    wire [15:0]out_mem_addr;
    wire [15:0]out_mem_addr_OBUF;
    wire out_mem_readEnable;
    wire out_mem_readEnable_OBUF;
    wire out_mem_readEnable_i_2_n_0;
    wire out_mem_writeEnable;
    wire out_mem_writeEnable_OBUF;
    wire out_mem_writeEnable_i_1_n_0;
    wire [12:0]p_1_in;
    wire [14:0]pc;
    wire pc[12]_i_3_n_0;
    wire pc[12]_i_4_n_0;
    wire pc[12]_i_5_n_0;
    wire pc[12]_i_6_n_0;
    wire pc[14]_i_1_n_0;
    wire pc[14]_i_3_n_0;
    wire pc[14]_i_5_n_0;
    wire pc[14]_i_6_n_0;
    wire pc[14]_i_7_n_0;
    wire pc[4]_i_3_n_0;
    wire pc[4]_i_4_n_0;
    wire pc[4]_i_5_n_0;
    wire pc[4]_i_6_n_0;
    wire pc[5]_i_2_n_0;
    wire pc[5]_i_3_n_0;
    wire pc[5]_i_4_n_0;
    wire pc[5]_i_5_n_0;
    wire pc[8]_i_3_n_0;
    wire pc[8]_i_4_n_0;
    wire pc[8]_i_5_n_0;
    wire pc[8]_i_6_n_0;
    wire pc[9]_i_2_n_0;
    wire pc[9]_i_3_n_0;
    wire pc[9]_i_4_n_0;
    wire pc_reg[12]_i_2_n_0;
    wire pc_reg[12]_i_2_n_1;
    wire pc_reg[12]_i_2_n_2;
    wire pc_reg[12]_i_2_n_3;
    wire pc_reg[14]_i_4_n_3;
    wire pc_reg[4]_i_2_n_0;
    wire pc_reg[4]_i_2_n_1;
    wire pc_reg[4]_i_2_n_2;
    wire pc_reg[4]_i_2_n_3;
    wire pc_reg[8]_i_2_n_0;
    wire pc_reg[8]_i_2_n_1;
    wire pc_reg[8]_i_2_n_2;
    wire pc_reg[8]_i_2_n_3;
    wire [14:2]sp;
    wire sp[10]_i_10_n_0;
    wire sp[10]_i_11_n_0;
    wire sp[10]_i_12_n_0;
    wire sp[10]_i_5_n_0;
    wire sp[10]_i_6_n_0;
    wire sp[10]_i_7_n_0;
    wire sp[10]_i_8_n_0;
    wire sp[10]_i_9_n_0;
    wire sp[14]_i_10_n_0;
    wire sp[14]_i_11_n_0;
    wire sp[14]_i_12_n_0;
    wire sp[14]_i_13_n_0;
    wire sp[14]_i_14_n_0;
    wire sp[14]_i_15_n_0;
    wire sp[14]_i_16_n_0;
    wire sp[14]_i_1_n_0;
    wire sp[14]_i_4_n_0;
    wire sp[14]_i_6_n_0;
    wire sp[14]_i_8_n_0;
    wire sp[14]_i_9_n_0;
    wire sp[2]_i_2_n_0;
    wire sp[6]_i_10_n_0;
    wire sp[6]_i_11_n_0;
    wire sp[6]_i_12_n_0;
    wire sp[6]_i_5_n_0;
    wire sp[6]_i_6_n_0;
    wire sp[6]_i_7_n_0;
    wire sp[6]_i_8_n_0;
    wire sp[6]_i_9_n_0;
    wire sp_reg[10]_i_3_n_0;
    wire sp_reg[10]_i_3_n_1;
    wire sp_reg[10]_i_3_n_2;
    wire sp_reg[10]_i_3_n_3;
    wire sp_reg[10]_i_3_n_4;
    wire sp_reg[10]_i_3_n_5;
    wire sp_reg[10]_i_3_n_6;
    wire sp_reg[10]_i_3_n_7;
    wire sp_reg[10]_i_4_n_0;
    wire sp_reg[10]_i_4_n_1;
    wire sp_reg[10]_i_4_n_2;
    wire sp_reg[10]_i_4_n_3;
    wire sp_reg[10]_i_4_n_4;
    wire sp_reg[10]_i_4_n_5;
    wire sp_reg[10]_i_4_n_6;
    wire sp_reg[10]_i_4_n_7;
    wire sp_reg[14]_i_5_n_1;
    wire sp_reg[14]_i_5_n_2;
    wire sp_reg[14]_i_5_n_3;
    wire sp_reg[14]_i_5_n_4;
    wire sp_reg[14]_i_5_n_5;
    wire sp_reg[14]_i_5_n_6;
    wire sp_reg[14]_i_5_n_7;
    wire sp_reg[14]_i_7_n_1;
    wire sp_reg[14]_i_7_n_2;
    wire sp_reg[14]_i_7_n_3;
    wire sp_reg[14]_i_7_n_4;
    wire sp_reg[14]_i_7_n_5;
    wire sp_reg[14]_i_7_n_6;
    wire sp_reg[14]_i_7_n_7;
    wire sp_reg[6]_i_3_n_0;
    wire sp_reg[6]_i_3_n_1;
    wire sp_reg[6]_i_3_n_2;
    wire sp_reg[6]_i_3_n_3;
    wire sp_reg[6]_i_3_n_4;
    wire sp_reg[6]_i_3_n_5;
    wire sp_reg[6]_i_3_n_6;
    wire sp_reg[6]_i_3_n_7;
    wire sp_reg[6]_i_4_n_0;
    wire sp_reg[6]_i_4_n_1;
    wire sp_reg[6]_i_4_n_2;
    wire sp_reg[6]_i_4_n_3;
    wire sp_reg[6]_i_4_n_4;
    wire sp_reg[6]_i_4_n_5;
    wire sp_reg[6]_i_4_n_6;
    wire sp_reg[6]_i_4_n_7;
    wire [14:2]sp_reg_n_0_;

    LUT6 FSM_sequential_state[0]_i_1
    (
        .O(FSM_sequential_state[0]_i_1_n_0),
        .I0(FSM_sequential_state[0]_i_2_n_0),
        .I1(FSM_sequential_state_reg_n_0_[2]),
        .I2(FSM_sequential_state[0]_i_3_n_0),
        .I3(FSM_sequential_state[0]_i_4_n_0),
        .I4(FSM_sequential_state[0]_i_5_n_0),
        .I5(FSM_sequential_state[0]_i_6_n_0)
    );
    LUT2 FSM_sequential_state[0]_i_2
    (
        .O(FSM_sequential_state[0]_i_2_n_0),
        .I0(FSM_sequential_state_reg_n_0_[0]),
        .I1(FSM_sequential_state_reg_n_0_[1])
    );
    LUT4 FSM_sequential_state[0]_i_3
    (
        .O(FSM_sequential_state[0]_i_3_n_0),
        .I0(FSM_sequential_state_reg_n_0_[3]),
        .I1(FSM_sequential_state_reg_n_0_[2]),
        .I2(FSM_sequential_state_reg_n_0_[1]),
        .I3(FSM_sequential_state_reg_n_0_[0])
    );
    LUT6 FSM_sequential_state[0]_i_4
    (
        .O(FSM_sequential_state[0]_i_4_n_0),
        .I0(decodedOpcode_reg_n_0_[2]),
        .I1(decodedOpcode_reg_n_0_[1]),
        .I2(decodedOpcode_reg_n_0_[0]),
        .I3(FSM_sequential_state_reg_n_0_[0]),
        .I4(in_mem_busy_IBUF),
        .I5(FSM_sequential_state_reg_n_0_[1])
    );
    LUT6 FSM_sequential_state[0]_i_5
    (
        .O(FSM_sequential_state[0]_i_5_n_0),
        .I0(FSM_sequential_state_reg_n_0_[0]),
        .I1(FSM_sequential_state_reg_n_0_[1]),
        .I2(decodedOpcode_reg_n_0_[2]),
        .I3(decodedOpcode_reg_n_0_[4]),
        .I4(decodedOpcode_reg_n_0_[3]),
        .I5(decodedOpcode_reg_n_0_[1])
    );
    LUT6 FSM_sequential_state[0]_i_6
    (
        .O(FSM_sequential_state[0]_i_6_n_0),
        .I0(in_mem_busy_IBUF),
        .I1(decodedOpcode_reg_n_0_[2]),
        .I2(decodedOpcode_reg_n_0_[3]),
        .I3(decodedOpcode_reg_n_0_[4]),
        .I4(FSM_sequential_state_reg_n_0_[1]),
        .I5(FSM_sequential_state_reg_n_0_[0])
    );
    LUT5 FSM_sequential_state[1]_i_3
    (
        .O(FSM_sequential_state[1]_i_3_n_0),
        .I0(FSM_sequential_state_reg_n_0_[2]),
        .I1(decodedOpcode_reg_n_0_[2]),
        .I2(decodedOpcode_reg_n_0_[4]),
        .I3(decodedOpcode_reg_n_0_[0]),
        .I4(decodedOpcode_reg_n_0_[3])
    );
    LUT5 FSM_sequential_state[2]_i_3
    (
        .O(FSM_sequential_state[2]_i_3_n_0),
        .I0(FSM_sequential_state_reg_n_0_[0]),
        .I1(FSM_sequential_state_reg_n_0_[1]),
        .I2(decodedOpcode_reg_n_0_[4]),
        .I3(decodedOpcode_reg_n_0_[3]),
        .I4(decodedOpcode_reg_n_0_[2])
    );
    LUT5 FSM_sequential_state[3]_i_1
    (
        .O(FSM_sequential_state[3]_i_1_n_0),
        .I0(FSM_sequential_state_reg_n_0_[3]),
        .I1(in_mem_busy_IBUF),
        .I2(FSM_sequential_state_reg_n_0_[0]),
        .I3(FSM_sequential_state_reg_n_0_[2]),
        .I4(FSM_sequential_state_reg_n_0_[1])
    );
    LUT4 FSM_sequential_state[3]_i_3
    (
        .O(FSM_sequential_state[3]_i_3_n_0),
        .I0(FSM_sequential_state_reg_n_0_[3]),
        .I1(FSM_sequential_state_reg_n_0_[0]),
        .I2(FSM_sequential_state_reg_n_0_[2]),
        .I3(FSM_sequential_state_reg_n_0_[1])
    );
    LUT5 FSM_sequential_state[3]_i_5
    (
        .O(FSM_sequential_state[3]_i_5_n_0),
        .I0(FSM_sequential_state_reg_n_0_[1]),
        .I1(FSM_sequential_state_reg_n_0_[0]),
        .I2(in_mem_busy_IBUF),
        .I3(FSM_sequential_state_reg_n_0_[3]),
        .I4(FSM_sequential_state_reg_n_0_[2])
    );
    FDCE FSM_sequential_state_reg[0]
    (
        .Q(FSM_sequential_state_reg_n_0_[0]),
        .C(clk_IBUF_BUFG),
        .CE(FSM_sequential_state[3]_i_1_n_0),
        .CLR(areset_IBUF),
        .D(FSM_sequential_state[0]_i_1_n_0)
    );
    FDCE FSM_sequential_state_reg[1]
    (
        .Q(FSM_sequential_state_reg_n_0_[1]),
        .C(clk_IBUF_BUFG),
        .CE(FSM_sequential_state[3]_i_1_n_0),
        .CLR(areset_IBUF),
        .D(memory_n_2)
    );
    FDCE FSM_sequential_state_reg[2]
    (
        .Q(FSM_sequential_state_reg_n_0_[2]),
        .C(clk_IBUF_BUFG),
        .CE(FSM_sequential_state[3]_i_1_n_0),
        .CLR(areset_IBUF),
        .D(memory_n_1)
    );
    FDCE FSM_sequential_state_reg[3]
    (
        .Q(FSM_sequential_state_reg_n_0_[3]),
        .C(clk_IBUF_BUFG),
        .CE(FSM_sequential_state[3]_i_1_n_0),
        .CLR(areset_IBUF),
        .D(memory_n_0)
    );
    GND GND
    (
        .G(<const0>)
    );
    VCC VCC
    (
        .P(<const1>)
    );
    IBUF areset_IBUF_inst
    (
        .O(areset_IBUF),
        .I(areset)
    );
    OBUF break_OBUF_inst
    (
        .O(break),
        .I(break_OBUF)
    );
    LUT6 break_i_1
    (
        .O(break_i_1_n_0),
        .I0(FSM_sequential_state[3]_i_3_n_0),
        .I1(decodedOpcode_reg_n_0_[0]),
        .I2(break_i_2_n_0),
        .I3(decodedOpcode_reg_n_0_[1]),
        .I4(decodedOpcode_reg_n_0_[4]),
        .I5(break_OBUF)
    );
    LUT2 break_i_2
    (
        .O(break_i_2_n_0),
        .I0(decodedOpcode_reg_n_0_[2]),
        .I1(decodedOpcode_reg_n_0_[3])
    );
    FDCE break_reg
    (
        .Q(break_OBUF),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(break_i_1_n_0)
    );
    BUFG clk_IBUF_BUFG_inst
    (
        .O(clk_IBUF_BUFG),
        .I(clk_IBUF)
    );
    IBUF clk_IBUF_inst
    (
        .O(clk_IBUF),
        .I(clk)
    );
    LUT4 decodedOpcode[4]_i_2
    (
        .O(decodedOpcode[4]_i_2_n_0),
        .I0(FSM_sequential_state_reg_n_0_[1]),
        .I1(FSM_sequential_state_reg_n_0_[3]),
        .I2(FSM_sequential_state_reg_n_0_[0]),
        .I3(FSM_sequential_state_reg_n_0_[2])
    );
    LUT3 decodedOpcode[4]_i_5
    (
        .O(decodedOpcode[4]_i_5_n_0),
        .I0(inInterrupt_reg_n_0),
        .I1(interrupt_IBUF),
        .I2(idim_flag)
    );
    FDRE decodedOpcode_reg[0]
    (
        .Q(decodedOpcode_reg_n_0_[0]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(decodedOpcode[0]),
        .R(<const0>)
    );
    FDRE decodedOpcode_reg[1]
    (
        .Q(decodedOpcode_reg_n_0_[1]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(decodedOpcode[1]),
        .R(<const0>)
    );
    FDRE decodedOpcode_reg[2]
    (
        .Q(decodedOpcode_reg_n_0_[2]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(decodedOpcode[2]),
        .R(<const0>)
    );
    FDRE decodedOpcode_reg[3]
    (
        .Q(decodedOpcode_reg_n_0_[3]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(decodedOpcode[3]),
        .R(<const0>)
    );
    FDRE decodedOpcode_reg[4]
    (
        .Q(decodedOpcode_reg_n_0_[4]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(decodedOpcode[4]),
        .R(<const0>)
    );
    LUT5 g0_b0
    (
        .O(g0_b0_n_0),
        .I0(decodedOpcode_reg_n_0_[0]),
        .I1(decodedOpcode_reg_n_0_[1]),
        .I2(decodedOpcode_reg_n_0_[2]),
        .I3(decodedOpcode_reg_n_0_[3]),
        .I4(decodedOpcode_reg_n_0_[4])
    );
    LUT5 g0_b0__0
    (
        .O(g0_b0__0_n_0),
        .I0(decodedOpcode_reg_n_0_[0]),
        .I1(decodedOpcode_reg_n_0_[1]),
        .I2(decodedOpcode_reg_n_0_[2]),
        .I3(decodedOpcode_reg_n_0_[3]),
        .I4(decodedOpcode_reg_n_0_[4])
    );
    LUT5 idim_flag_i_1
    (
        .O(idim_flag_i_1_n_0),
        .I0(decodedOpcode_reg_n_0_[3]),
        .I1(decodedOpcode_reg_n_0_[4]),
        .I2(decodedOpcode_reg_n_0_[1]),
        .I3(decodedOpcode_reg_n_0_[2]),
        .I4(decodedOpcode_reg_n_0_[0])
    );
    FDCE idim_flag_reg
    (
        .Q(idim_flag),
        .C(clk_IBUF_BUFG),
        .CE(pc[14]_i_1_n_0),
        .CLR(areset_IBUF),
        .D(idim_flag_i_1_n_0)
    );
    LUT4 inInterrupt_i_1
    (
        .O(inInterrupt_i_1_n_0),
        .I0(decodedOpcode[4]_i_2_n_0),
        .I1(idim_flag),
        .I2(inInterrupt_reg_n_0),
        .I3(interrupt_IBUF)
    );
    FDCE inInterrupt_reg
    (
        .Q(inInterrupt_reg_n_0),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(inInterrupt_i_1_n_0)
    );
    IBUF in_mem_busy_IBUF_inst
    (
        .O(in_mem_busy_IBUF),
        .I(in_mem_busy)
    );
    IBUF interrupt_IBUF_inst
    (
        .O(interrupt_IBUF),
        .I(interrupt)
    );
    LUT4 memAAddr[10]_i_4
    (
        .O(memAAddr[10]_i_4_n_0),
        .I0(decodedOpcode_reg_n_0_[2]),
        .I1(decodedOpcode_reg_n_0_[0]),
        .I2(decodedOpcode_reg_n_0_[1]),
        .I3(memBAddr_reg[13]_i_2_n_7)
    );
    LUT4 memAAddr[11]_i_4
    (
        .O(memAAddr[11]_i_4_n_0),
        .I0(decodedOpcode_reg_n_0_[2]),
        .I1(decodedOpcode_reg_n_0_[0]),
        .I2(decodedOpcode_reg_n_0_[1]),
        .I3(memBAddr_reg[13]_i_2_n_6)
    );
    LUT4 memAAddr[12]_i_4
    (
        .O(memAAddr[12]_i_4_n_0),
        .I0(decodedOpcode_reg_n_0_[2]),
        .I1(decodedOpcode_reg_n_0_[0]),
        .I2(decodedOpcode_reg_n_0_[1]),
        .I3(memBAddr_reg[13]_i_2_n_5)
    );
    LUT4 memAAddr[13]_i_4
    (
        .O(memAAddr[13]_i_4_n_0),
        .I0(decodedOpcode_reg_n_0_[2]),
        .I1(decodedOpcode_reg_n_0_[0]),
        .I2(decodedOpcode_reg_n_0_[1]),
        .I3(memBAddr_reg[13]_i_2_n_4)
    );
    LUT6 memAAddr[14]_i_4
    (
        .O(memAAddr[14]_i_4_n_0),
        .I0(decodedOpcode_reg_n_0_[4]),
        .I1(decodedOpcode_reg_n_0_[3]),
        .I2(decodedOpcode_reg_n_0_[2]),
        .I3(decodedOpcode_reg_n_0_[0]),
        .I4(idim_flag),
        .I5(decodedOpcode_reg_n_0_[1])
    );
    LUT6 memAAddr[14]_i_5
    (
        .O(memAAddr[14]_i_5_n_0),
        .I0(decodedOpcode_reg_n_0_[1]),
        .I1(idim_flag),
        .I2(decodedOpcode_reg_n_0_[4]),
        .I3(decodedOpcode_reg_n_0_[2]),
        .I4(decodedOpcode_reg_n_0_[3]),
        .I5(decodedOpcode_reg_n_0_[0])
    );
    LUT4 memAAddr[14]_i_6
    (
        .O(memAAddr[14]_i_6_n_0),
        .I0(decodedOpcode_reg_n_0_[2]),
        .I1(decodedOpcode_reg_n_0_[0]),
        .I2(decodedOpcode_reg_n_0_[1]),
        .I3(memBAddr_reg[14]_i_2_n_7)
    );
    LUT4 memAAddr[2]_i_3
    (
        .O(memAAddr[2]_i_3_n_0),
        .I0(decodedOpcode_reg_n_0_[0]),
        .I1(decodedOpcode_reg_n_0_[3]),
        .I2(decodedOpcode_reg_n_0_[2]),
        .I3(decodedOpcode_reg_n_0_[1])
    );
    LUT4 memAAddr[2]_i_4
    (
        .O(memAAddr[2]_i_4_n_0),
        .I0(decodedOpcode_reg_n_0_[2]),
        .I1(decodedOpcode_reg_n_0_[0]),
        .I2(decodedOpcode_reg_n_0_[1]),
        .I3(memBAddr_reg[5]_i_2_n_7)
    );
    LUT4 memAAddr[3]_i_4
    (
        .O(memAAddr[3]_i_4_n_0),
        .I0(decodedOpcode_reg_n_0_[2]),
        .I1(decodedOpcode_reg_n_0_[0]),
        .I2(decodedOpcode_reg_n_0_[1]),
        .I3(memBAddr_reg[5]_i_2_n_6)
    );
    LUT4 memAAddr[4]_i_4
    (
        .O(memAAddr[4]_i_4_n_0),
        .I0(decodedOpcode_reg_n_0_[2]),
        .I1(decodedOpcode_reg_n_0_[0]),
        .I2(decodedOpcode_reg_n_0_[1]),
        .I3(memBAddr_reg[5]_i_2_n_5)
    );
    LUT4 memAAddr[5]_i_4
    (
        .O(memAAddr[5]_i_4_n_0),
        .I0(decodedOpcode_reg_n_0_[2]),
        .I1(decodedOpcode_reg_n_0_[0]),
        .I2(decodedOpcode_reg_n_0_[1]),
        .I3(memBAddr_reg[5]_i_2_n_4)
    );
    LUT4 memAAddr[6]_i_4
    (
        .O(memAAddr[6]_i_4_n_0),
        .I0(decodedOpcode_reg_n_0_[2]),
        .I1(decodedOpcode_reg_n_0_[0]),
        .I2(decodedOpcode_reg_n_0_[1]),
        .I3(memBAddr_reg[9]_i_2_n_7)
    );
    LUT4 memAAddr[7]_i_4
    (
        .O(memAAddr[7]_i_4_n_0),
        .I0(decodedOpcode_reg_n_0_[2]),
        .I1(decodedOpcode_reg_n_0_[0]),
        .I2(decodedOpcode_reg_n_0_[1]),
        .I3(memBAddr_reg[9]_i_2_n_6)
    );
    LUT4 memAAddr[8]_i_4
    (
        .O(memAAddr[8]_i_4_n_0),
        .I0(decodedOpcode_reg_n_0_[2]),
        .I1(decodedOpcode_reg_n_0_[0]),
        .I2(decodedOpcode_reg_n_0_[1]),
        .I3(memBAddr_reg[9]_i_2_n_5)
    );
    LUT4 memAAddr[9]_i_4
    (
        .O(memAAddr[9]_i_4_n_0),
        .I0(decodedOpcode_reg_n_0_[2]),
        .I1(decodedOpcode_reg_n_0_[0]),
        .I2(decodedOpcode_reg_n_0_[1]),
        .I3(memBAddr_reg[9]_i_2_n_4)
    );
    FDCE memAAddr_reg[10]
    (
        .Q(memAAddr_reg_n_0_[10]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memAAddr[10])
    );
    FDCE memAAddr_reg[11]
    (
        .Q(memAAddr_reg_n_0_[11]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memAAddr[11])
    );
    FDCE memAAddr_reg[12]
    (
        .Q(memAAddr_reg_n_0_[12]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memAAddr[12])
    );
    FDCE memAAddr_reg[13]
    (
        .Q(memAAddr_reg_n_0_[13]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memAAddr[13])
    );
    FDCE memAAddr_reg[14]
    (
        .Q(memAAddr_reg_n_0_[14]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memAAddr[14])
    );
    FDCE memAAddr_reg[2]
    (
        .Q(memAAddr_reg_n_0_[2]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memAAddr[2])
    );
    FDCE memAAddr_reg[3]
    (
        .Q(memAAddr_reg_n_0_[3]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memAAddr[3])
    );
    FDCE memAAddr_reg[4]
    (
        .Q(memAAddr_reg_n_0_[4]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memAAddr[4])
    );
    FDCE memAAddr_reg[5]
    (
        .Q(memAAddr_reg_n_0_[5]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memAAddr[5])
    );
    FDCE memAAddr_reg[6]
    (
        .Q(memAAddr_reg_n_0_[6]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memAAddr[6])
    );
    FDCE memAAddr_reg[7]
    (
        .Q(memAAddr_reg_n_0_[7]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memAAddr[7])
    );
    FDCE memAAddr_reg[8]
    (
        .Q(memAAddr_reg_n_0_[8]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memAAddr[8])
    );
    FDCE memAAddr_reg[9]
    (
        .Q(memAAddr_reg_n_0_[9]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memAAddr[9])
    );
    LUT6 memAWriteEnable_i_1
    (
        .O(memAWriteEnable),
        .I0(g0_b0_n_0),
        .I1(FSM_sequential_state_reg_n_0_[1]),
        .I2(in_mem_busy_IBUF),
        .I3(FSM_sequential_state_reg_n_0_[2]),
        .I4(FSM_sequential_state_reg_n_0_[0]),
        .I5(FSM_sequential_state_reg_n_0_[3])
    );
    FDCE memAWriteEnable_reg
    (
        .Q(memAWriteEnable_reg_n_0),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memAWriteEnable)
    );
    LUT5 memAWrite[0]_i_4
    (
        .O(memAWrite[0]_i_4_n_0),
        .I0(opcode_reg_n_0_[0]),
        .I1(data0[0]),
        .I2(decodedOpcode_reg_n_0_[1]),
        .I3(decodedOpcode_reg_n_0_[0]),
        .I4(decodedOpcode_reg_n_0_[2])
    );
    LUT5 memAWrite[10]_i_4
    (
        .O(memAWrite[10]_i_4_n_0),
        .I0(p_1_in[8]),
        .I1(decodedOpcode_reg_n_0_[0]),
        .I2(decodedOpcode_reg_n_0_[2]),
        .I3(decodedOpcode_reg_n_0_[1]),
        .I4(sp_reg_n_0_[10])
    );
    LUT6 memAWrite[10]_i_7
    (
        .O(memAWrite[10]_i_7_n_0),
        .I0(data2[10]),
        .I1(decodedOpcode_reg_n_0_[3]),
        .I2(idim_flag),
        .I3(opcode_reg_n_0_[6]),
        .I4(decodedOpcode_reg_n_0_[0]),
        .I5(decodedOpcode_reg_n_0_[2])
    );
    LUT5 memAWrite[11]_i_4
    (
        .O(memAWrite[11]_i_4_n_0),
        .I0(p_1_in[9]),
        .I1(decodedOpcode_reg_n_0_[0]),
        .I2(decodedOpcode_reg_n_0_[2]),
        .I3(decodedOpcode_reg_n_0_[1]),
        .I4(sp_reg_n_0_[11])
    );
    LUT6 memAWrite[11]_i_7
    (
        .O(memAWrite[11]_i_7_n_0),
        .I0(data2[11]),
        .I1(decodedOpcode_reg_n_0_[3]),
        .I2(idim_flag),
        .I3(opcode_reg_n_0_[6]),
        .I4(decodedOpcode_reg_n_0_[0]),
        .I5(decodedOpcode_reg_n_0_[2])
    );
    LUT5 memAWrite[12]_i_4
    (
        .O(memAWrite[12]_i_4_n_0),
        .I0(p_1_in[10]),
        .I1(decodedOpcode_reg_n_0_[0]),
        .I2(decodedOpcode_reg_n_0_[2]),
        .I3(decodedOpcode_reg_n_0_[1]),
        .I4(sp_reg_n_0_[12])
    );
    LUT6 memAWrite[12]_i_7
    (
        .O(memAWrite[12]_i_7_n_0),
        .I0(data2[12]),
        .I1(decodedOpcode_reg_n_0_[3]),
        .I2(idim_flag),
        .I3(opcode_reg_n_0_[6]),
        .I4(decodedOpcode_reg_n_0_[0]),
        .I5(decodedOpcode_reg_n_0_[2])
    );
    LUT5 memAWrite[13]_i_4
    (
        .O(memAWrite[13]_i_4_n_0),
        .I0(p_1_in[11]),
        .I1(decodedOpcode_reg_n_0_[0]),
        .I2(decodedOpcode_reg_n_0_[2]),
        .I3(decodedOpcode_reg_n_0_[1]),
        .I4(sp_reg_n_0_[13])
    );
    LUT6 memAWrite[13]_i_7
    (
        .O(memAWrite[13]_i_7_n_0),
        .I0(data2[13]),
        .I1(decodedOpcode_reg_n_0_[3]),
        .I2(idim_flag),
        .I3(opcode_reg_n_0_[6]),
        .I4(decodedOpcode_reg_n_0_[0]),
        .I5(decodedOpcode_reg_n_0_[2])
    );
    LUT5 memAWrite[14]_i_4
    (
        .O(memAWrite[14]_i_4_n_0),
        .I0(p_1_in[12]),
        .I1(decodedOpcode_reg_n_0_[0]),
        .I2(decodedOpcode_reg_n_0_[2]),
        .I3(decodedOpcode_reg_n_0_[1]),
        .I4(sp_reg_n_0_[14])
    );
    LUT6 memAWrite[14]_i_7
    (
        .O(memAWrite[14]_i_7_n_0),
        .I0(data2[14]),
        .I1(decodedOpcode_reg_n_0_[3]),
        .I2(idim_flag),
        .I3(opcode_reg_n_0_[6]),
        .I4(decodedOpcode_reg_n_0_[0]),
        .I5(decodedOpcode_reg_n_0_[2])
    );
    LUT5 memAWrite[1]_i_4
    (
        .O(memAWrite[1]_i_4_n_0),
        .I0(opcode_reg_n_0_[1]),
        .I1(data0[1]),
        .I2(decodedOpcode_reg_n_0_[1]),
        .I3(decodedOpcode_reg_n_0_[0]),
        .I4(decodedOpcode_reg_n_0_[2])
    );
    LUT5 memAWrite[2]_i_4
    (
        .O(memAWrite[2]_i_4_n_0),
        .I0(p_1_in[0]),
        .I1(decodedOpcode_reg_n_0_[0]),
        .I2(decodedOpcode_reg_n_0_[2]),
        .I3(decodedOpcode_reg_n_0_[1]),
        .I4(sp_reg_n_0_[2])
    );
    LUT5 memAWrite[2]_i_5
    (
        .O(memAWrite[2]_i_5_n_0),
        .I0(data2[2]),
        .I1(decodedOpcode_reg_n_0_[3]),
        .I2(opcode_reg_n_0_[2]),
        .I3(decodedOpcode_reg_n_0_[0]),
        .I4(decodedOpcode_reg_n_0_[2])
    );
    LUT3 memAWrite[31]_i_4
    (
        .O(memAWrite[31]_i_4_n_0),
        .I0(decodedOpcode_reg_n_0_[2]),
        .I1(decodedOpcode_reg_n_0_[3]),
        .I2(decodedOpcode_reg_n_0_[0])
    );
    LUT5 memAWrite[3]_i_4
    (
        .O(memAWrite[3]_i_4_n_0),
        .I0(p_1_in[1]),
        .I1(decodedOpcode_reg_n_0_[0]),
        .I2(decodedOpcode_reg_n_0_[2]),
        .I3(decodedOpcode_reg_n_0_[1]),
        .I4(sp_reg_n_0_[3])
    );
    LUT5 memAWrite[3]_i_5
    (
        .O(memAWrite[3]_i_5_n_0),
        .I0(data2[3]),
        .I1(decodedOpcode_reg_n_0_[3]),
        .I2(opcode_reg_n_0_[3]),
        .I3(decodedOpcode_reg_n_0_[0]),
        .I4(decodedOpcode_reg_n_0_[2])
    );
    LUT5 memAWrite[4]_i_4
    (
        .O(memAWrite[4]_i_4_n_0),
        .I0(p_1_in[2]),
        .I1(decodedOpcode_reg_n_0_[0]),
        .I2(decodedOpcode_reg_n_0_[2]),
        .I3(decodedOpcode_reg_n_0_[1]),
        .I4(sp_reg_n_0_[4])
    );
    LUT5 memAWrite[4]_i_5
    (
        .O(memAWrite[4]_i_5_n_0),
        .I0(data2[4]),
        .I1(decodedOpcode_reg_n_0_[3]),
        .I2(opcode_reg_n_0_[4]),
        .I3(decodedOpcode_reg_n_0_[0]),
        .I4(decodedOpcode_reg_n_0_[2])
    );
    LUT5 memAWrite[5]_i_4
    (
        .O(memAWrite[5]_i_4_n_0),
        .I0(p_1_in[3]),
        .I1(decodedOpcode_reg_n_0_[0]),
        .I2(decodedOpcode_reg_n_0_[2]),
        .I3(decodedOpcode_reg_n_0_[1]),
        .I4(sp_reg_n_0_[5])
    );
    LUT5 memAWrite[5]_i_5
    (
        .O(memAWrite[5]_i_5_n_0),
        .I0(data2[5]),
        .I1(decodedOpcode_reg_n_0_[3]),
        .I2(opcode_reg_n_0_[5]),
        .I3(decodedOpcode_reg_n_0_[0]),
        .I4(decodedOpcode_reg_n_0_[2])
    );
    LUT5 memAWrite[6]_i_4
    (
        .O(memAWrite[6]_i_4_n_0),
        .I0(p_1_in[4]),
        .I1(decodedOpcode_reg_n_0_[0]),
        .I2(decodedOpcode_reg_n_0_[2]),
        .I3(decodedOpcode_reg_n_0_[1]),
        .I4(sp_reg_n_0_[6])
    );
    LUT5 memAWrite[6]_i_5
    (
        .O(memAWrite[6]_i_5_n_0),
        .I0(data2[6]),
        .I1(decodedOpcode_reg_n_0_[3]),
        .I2(opcode_reg_n_0_[6]),
        .I3(decodedOpcode_reg_n_0_[0]),
        .I4(decodedOpcode_reg_n_0_[2])
    );
    LUT5 memAWrite[7]_i_4
    (
        .O(memAWrite[7]_i_4_n_0),
        .I0(p_1_in[5]),
        .I1(decodedOpcode_reg_n_0_[0]),
        .I2(decodedOpcode_reg_n_0_[2]),
        .I3(decodedOpcode_reg_n_0_[1]),
        .I4(sp_reg_n_0_[7])
    );
    LUT6 memAWrite[7]_i_7
    (
        .O(memAWrite[7]_i_7_n_0),
        .I0(data2[7]),
        .I1(decodedOpcode_reg_n_0_[3]),
        .I2(idim_flag),
        .I3(opcode_reg_n_0_[6]),
        .I4(decodedOpcode_reg_n_0_[0]),
        .I5(decodedOpcode_reg_n_0_[2])
    );
    LUT5 memAWrite[8]_i_4
    (
        .O(memAWrite[8]_i_4_n_0),
        .I0(p_1_in[6]),
        .I1(decodedOpcode_reg_n_0_[0]),
        .I2(decodedOpcode_reg_n_0_[2]),
        .I3(decodedOpcode_reg_n_0_[1]),
        .I4(sp_reg_n_0_[8])
    );
    LUT6 memAWrite[8]_i_7
    (
        .O(memAWrite[8]_i_7_n_0),
        .I0(data2[8]),
        .I1(decodedOpcode_reg_n_0_[3]),
        .I2(idim_flag),
        .I3(opcode_reg_n_0_[6]),
        .I4(decodedOpcode_reg_n_0_[0]),
        .I5(decodedOpcode_reg_n_0_[2])
    );
    LUT5 memAWrite[9]_i_4
    (
        .O(memAWrite[9]_i_4_n_0),
        .I0(p_1_in[7]),
        .I1(decodedOpcode_reg_n_0_[0]),
        .I2(decodedOpcode_reg_n_0_[2]),
        .I3(decodedOpcode_reg_n_0_[1]),
        .I4(sp_reg_n_0_[9])
    );
    LUT6 memAWrite[9]_i_7
    (
        .O(memAWrite[9]_i_7_n_0),
        .I0(data2[9]),
        .I1(decodedOpcode_reg_n_0_[3]),
        .I2(idim_flag),
        .I3(opcode_reg_n_0_[6]),
        .I4(decodedOpcode_reg_n_0_[0]),
        .I5(decodedOpcode_reg_n_0_[2])
    );
    FDCE memAWrite_reg[0]
    (
        .Q(memAWrite_reg_n_0_[0]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memAWrite[0])
    );
    FDCE memAWrite_reg[10]
    (
        .Q(memAWrite_reg_n_0_[10]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memAWrite[10])
    );
    FDCE memAWrite_reg[11]
    (
        .Q(memAWrite_reg_n_0_[11]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memAWrite[11])
    );
    FDCE memAWrite_reg[12]
    (
        .Q(memAWrite_reg_n_0_[12]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memAWrite[12])
    );
    FDCE memAWrite_reg[13]
    (
        .Q(memAWrite_reg_n_0_[13]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memAWrite[13])
    );
    FDCE memAWrite_reg[14]
    (
        .Q(memAWrite_reg_n_0_[14]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memAWrite[14])
    );
    FDCE memAWrite_reg[15]
    (
        .Q(memAWrite_reg_n_0_[15]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memAWrite[15])
    );
    FDCE memAWrite_reg[16]
    (
        .Q(memAWrite_reg_n_0_[16]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memAWrite[16])
    );
    FDCE memAWrite_reg[17]
    (
        .Q(memAWrite_reg_n_0_[17]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memAWrite[17])
    );
    FDCE memAWrite_reg[18]
    (
        .Q(memAWrite_reg_n_0_[18]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memAWrite[18])
    );
    FDCE memAWrite_reg[19]
    (
        .Q(memAWrite_reg_n_0_[19]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memAWrite[19])
    );
    FDCE memAWrite_reg[1]
    (
        .Q(memAWrite_reg_n_0_[1]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memAWrite[1])
    );
    FDCE memAWrite_reg[20]
    (
        .Q(memAWrite_reg_n_0_[20]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memAWrite[20])
    );
    FDCE memAWrite_reg[21]
    (
        .Q(memAWrite_reg_n_0_[21]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memAWrite[21])
    );
    FDCE memAWrite_reg[22]
    (
        .Q(memAWrite_reg_n_0_[22]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memAWrite[22])
    );
    FDCE memAWrite_reg[23]
    (
        .Q(memAWrite_reg_n_0_[23]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memAWrite[23])
    );
    FDCE memAWrite_reg[24]
    (
        .Q(memAWrite_reg_n_0_[24]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memAWrite[24])
    );
    FDCE memAWrite_reg[25]
    (
        .Q(memAWrite_reg_n_0_[25]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memAWrite[25])
    );
    FDCE memAWrite_reg[26]
    (
        .Q(memAWrite_reg_n_0_[26]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memAWrite[26])
    );
    FDCE memAWrite_reg[27]
    (
        .Q(memAWrite_reg_n_0_[27]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memAWrite[27])
    );
    FDCE memAWrite_reg[28]
    (
        .Q(memAWrite_reg_n_0_[28]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memAWrite[28])
    );
    FDCE memAWrite_reg[29]
    (
        .Q(memAWrite_reg_n_0_[29]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memAWrite[29])
    );
    FDCE memAWrite_reg[2]
    (
        .Q(memAWrite_reg_n_0_[2]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memAWrite[2])
    );
    FDCE memAWrite_reg[30]
    (
        .Q(memAWrite_reg_n_0_[30]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memAWrite[30])
    );
    FDCE memAWrite_reg[31]
    (
        .Q(memAWrite_reg_n_0_[31]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memAWrite[31])
    );
    FDCE memAWrite_reg[3]
    (
        .Q(memAWrite_reg_n_0_[3]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memAWrite[3])
    );
    FDCE memAWrite_reg[4]
    (
        .Q(memAWrite_reg_n_0_[4]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memAWrite[4])
    );
    FDCE memAWrite_reg[5]
    (
        .Q(memAWrite_reg_n_0_[5]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memAWrite[5])
    );
    FDCE memAWrite_reg[6]
    (
        .Q(memAWrite_reg_n_0_[6]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memAWrite[6])
    );
    FDCE memAWrite_reg[7]
    (
        .Q(memAWrite_reg_n_0_[7]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memAWrite[7])
    );
    FDCE memAWrite_reg[8]
    (
        .Q(memAWrite_reg_n_0_[8]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memAWrite[8])
    );
    FDCE memAWrite_reg[9]
    (
        .Q(memAWrite_reg_n_0_[9]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memAWrite[9])
    );
    LUT6 memBAddr[10]_i_1
    (
        .O(memBAddr[10]),
        .I0(FSM_sequential_state_reg_n_0_[1]),
        .I1(sp_reg[10]_i_3_n_4),
        .I2(decodedOpcode_reg_n_0_[4]),
        .I3(memBAddr_reg[13]_i_2_n_7),
        .I4(FSM_sequential_state_reg_n_0_[2]),
        .I5(p_1_in[8])
    );
    LUT6 memBAddr[11]_i_1
    (
        .O(memBAddr[11]),
        .I0(FSM_sequential_state_reg_n_0_[1]),
        .I1(sp_reg[14]_i_5_n_7),
        .I2(decodedOpcode_reg_n_0_[4]),
        .I3(memBAddr_reg[13]_i_2_n_6),
        .I4(FSM_sequential_state_reg_n_0_[2]),
        .I5(p_1_in[9])
    );
    LUT6 memBAddr[12]_i_1
    (
        .O(memBAddr[12]),
        .I0(FSM_sequential_state_reg_n_0_[1]),
        .I1(sp_reg[14]_i_5_n_6),
        .I2(decodedOpcode_reg_n_0_[4]),
        .I3(memBAddr_reg[13]_i_2_n_5),
        .I4(FSM_sequential_state_reg_n_0_[2]),
        .I5(p_1_in[10])
    );
    LUT6 memBAddr[13]_i_1
    (
        .O(memBAddr[13]),
        .I0(FSM_sequential_state_reg_n_0_[1]),
        .I1(sp_reg[14]_i_5_n_5),
        .I2(decodedOpcode_reg_n_0_[4]),
        .I3(memBAddr_reg[13]_i_2_n_4),
        .I4(FSM_sequential_state_reg_n_0_[2]),
        .I5(p_1_in[11])
    );
    LUT1 memBAddr[13]_i_3
    (
        .O(memBAddr[13]_i_3_n_0),
        .I0(sp_reg_n_0_[13])
    );
    LUT1 memBAddr[13]_i_4
    (
        .O(memBAddr[13]_i_4_n_0),
        .I0(sp_reg_n_0_[12])
    );
    LUT1 memBAddr[13]_i_5
    (
        .O(memBAddr[13]_i_5_n_0),
        .I0(sp_reg_n_0_[11])
    );
    LUT1 memBAddr[13]_i_6
    (
        .O(memBAddr[13]_i_6_n_0),
        .I0(sp_reg_n_0_[10])
    );
    LUT6 memBAddr[14]_i_1
    (
        .O(memBAddr[14]),
        .I0(FSM_sequential_state_reg_n_0_[1]),
        .I1(sp_reg[14]_i_5_n_4),
        .I2(decodedOpcode_reg_n_0_[4]),
        .I3(memBAddr_reg[14]_i_2_n_7),
        .I4(FSM_sequential_state_reg_n_0_[2]),
        .I5(p_1_in[12])
    );
    LUT1 memBAddr[14]_i_3
    (
        .O(memBAddr[14]_i_3_n_0),
        .I0(sp_reg_n_0_[14])
    );
    LUT6 memBAddr[2]_i_1
    (
        .O(memBAddr[2]),
        .I0(FSM_sequential_state_reg_n_0_[1]),
        .I1(sp_reg_n_0_[2]),
        .I2(decodedOpcode_reg_n_0_[4]),
        .I3(memBAddr_reg[5]_i_2_n_7),
        .I4(FSM_sequential_state_reg_n_0_[2]),
        .I5(p_1_in[0])
    );
    LUT6 memBAddr[3]_i_1
    (
        .O(memBAddr[3]),
        .I0(FSM_sequential_state_reg_n_0_[1]),
        .I1(sp_reg[6]_i_3_n_7),
        .I2(decodedOpcode_reg_n_0_[4]),
        .I3(memBAddr_reg[5]_i_2_n_6),
        .I4(FSM_sequential_state_reg_n_0_[2]),
        .I5(p_1_in[1])
    );
    LUT6 memBAddr[4]_i_1
    (
        .O(memBAddr[4]),
        .I0(FSM_sequential_state_reg_n_0_[1]),
        .I1(sp_reg[6]_i_3_n_6),
        .I2(decodedOpcode_reg_n_0_[4]),
        .I3(memBAddr_reg[5]_i_2_n_5),
        .I4(FSM_sequential_state_reg_n_0_[2]),
        .I5(p_1_in[2])
    );
    LUT6 memBAddr[5]_i_1
    (
        .O(memBAddr[5]),
        .I0(FSM_sequential_state_reg_n_0_[1]),
        .I1(sp_reg[6]_i_3_n_5),
        .I2(decodedOpcode_reg_n_0_[4]),
        .I3(memBAddr_reg[5]_i_2_n_4),
        .I4(FSM_sequential_state_reg_n_0_[2]),
        .I5(p_1_in[3])
    );
    LUT2 memBAddr[5]_i_3
    (
        .O(memBAddr[5]_i_3_n_0),
        .I0(sp_reg_n_0_[5]),
        .I1(opcode_reg_n_0_[3])
    );
    LUT2 memBAddr[5]_i_4
    (
        .O(memBAddr[5]_i_4_n_0),
        .I0(sp_reg_n_0_[4]),
        .I1(opcode_reg_n_0_[2])
    );
    LUT2 memBAddr[5]_i_5
    (
        .O(memBAddr[5]_i_5_n_0),
        .I0(sp_reg_n_0_[3]),
        .I1(opcode_reg_n_0_[1])
    );
    LUT2 memBAddr[5]_i_6
    (
        .O(memBAddr[5]_i_6_n_0),
        .I0(sp_reg_n_0_[2]),
        .I1(opcode_reg_n_0_[0])
    );
    LUT6 memBAddr[6]_i_1
    (
        .O(memBAddr[6]),
        .I0(FSM_sequential_state_reg_n_0_[1]),
        .I1(sp_reg[6]_i_3_n_4),
        .I2(decodedOpcode_reg_n_0_[4]),
        .I3(memBAddr_reg[9]_i_2_n_7),
        .I4(FSM_sequential_state_reg_n_0_[2]),
        .I5(p_1_in[4])
    );
    LUT6 memBAddr[7]_i_1
    (
        .O(memBAddr[7]),
        .I0(FSM_sequential_state_reg_n_0_[1]),
        .I1(sp_reg[10]_i_3_n_7),
        .I2(decodedOpcode_reg_n_0_[4]),
        .I3(memBAddr_reg[9]_i_2_n_6),
        .I4(FSM_sequential_state_reg_n_0_[2]),
        .I5(p_1_in[5])
    );
    LUT6 memBAddr[8]_i_1
    (
        .O(memBAddr[8]),
        .I0(FSM_sequential_state_reg_n_0_[1]),
        .I1(sp_reg[10]_i_3_n_6),
        .I2(decodedOpcode_reg_n_0_[4]),
        .I3(memBAddr_reg[9]_i_2_n_5),
        .I4(FSM_sequential_state_reg_n_0_[2]),
        .I5(p_1_in[6])
    );
    LUT6 memBAddr[9]_i_1
    (
        .O(memBAddr[9]),
        .I0(FSM_sequential_state_reg_n_0_[1]),
        .I1(sp_reg[10]_i_3_n_5),
        .I2(decodedOpcode_reg_n_0_[4]),
        .I3(memBAddr_reg[9]_i_2_n_4),
        .I4(FSM_sequential_state_reg_n_0_[2]),
        .I5(p_1_in[7])
    );
    LUT1 memBAddr[9]_i_3
    (
        .O(memBAddr[9]_i_3_n_0),
        .I0(sp_reg_n_0_[9])
    );
    LUT1 memBAddr[9]_i_4
    (
        .O(memBAddr[9]_i_4_n_0),
        .I0(sp_reg_n_0_[8])
    );
    LUT1 memBAddr[9]_i_5
    (
        .O(memBAddr[9]_i_5_n_0),
        .I0(sp_reg_n_0_[7])
    );
    LUT2 memBAddr[9]_i_6
    (
        .O(memBAddr[9]_i_6_n_0),
        .I0(sp_reg_n_0_[6]),
        .I1(opcode_reg_n_0_[4])
    );
    FDCE memBAddr_reg[10]
    (
        .Q(memBAddr_reg_n_0_[10]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memBAddr[10])
    );
    FDCE memBAddr_reg[11]
    (
        .Q(memBAddr_reg_n_0_[11]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memBAddr[11])
    );
    FDCE memBAddr_reg[12]
    (
        .Q(memBAddr_reg_n_0_[12]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memBAddr[12])
    );
    FDCE memBAddr_reg[13]
    (
        .Q(memBAddr_reg_n_0_[13]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memBAddr[13])
    );
    CARRY4 memBAddr_reg[13]_i_2
    (
        .CI(memBAddr_reg[9]_i_2_n_0),
        .CYINIT(<const0>),
        .CO[3:0]({memBAddr_reg[13]_i_2_n_0, memBAddr_reg[13]_i_2_n_1, memBAddr_reg[13]_i_2_n_2, memBAddr_reg[13]_i_2_n_3}),
        .O[3:0]({memBAddr_reg[13]_i_2_n_4, memBAddr_reg[13]_i_2_n_5, memBAddr_reg[13]_i_2_n_6, memBAddr_reg[13]_i_2_n_7}),
        .DI[3:0]({<const0>, <const0>, <const0>, <const0>}),
        .S[3:0]({memBAddr[13]_i_3_n_0, memBAddr[13]_i_4_n_0, memBAddr[13]_i_5_n_0, memBAddr[13]_i_6_n_0})
    );
    FDCE memBAddr_reg[14]
    (
        .Q(memBAddr_reg_n_0_[14]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memBAddr[14])
    );
    CARRY4 memBAddr_reg[14]_i_2
    (
        .CI(memBAddr_reg[13]_i_2_n_0),
        .CYINIT(<const0>),
        .CO[3:0](),
        .O[3:0]({}),
        .DI[3:0]({<const0>, <const0>, <const0>, <const0>}),
        .S[3:0]({<const0>, <const0>, <const0>, memBAddr[14]_i_3_n_0})
    );
    FDCE memBAddr_reg[2]
    (
        .Q(memBAddr_reg_n_0_[2]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memBAddr[2])
    );
    FDCE memBAddr_reg[3]
    (
        .Q(memBAddr_reg_n_0_[3]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memBAddr[3])
    );
    FDCE memBAddr_reg[4]
    (
        .Q(memBAddr_reg_n_0_[4]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memBAddr[4])
    );
    FDCE memBAddr_reg[5]
    (
        .Q(memBAddr_reg_n_0_[5]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memBAddr[5])
    );
    CARRY4 memBAddr_reg[5]_i_2
    (
        .CI(<const0>),
        .CYINIT(<const0>),
        .CO[3:0]({memBAddr_reg[5]_i_2_n_0, memBAddr_reg[5]_i_2_n_1, memBAddr_reg[5]_i_2_n_2, memBAddr_reg[5]_i_2_n_3}),
        .O[3:0]({memBAddr_reg[5]_i_2_n_4, memBAddr_reg[5]_i_2_n_5, memBAddr_reg[5]_i_2_n_6, memBAddr_reg[5]_i_2_n_7}),
        .DI[3:0]({sp_reg_n_0_[5], sp_reg_n_0_[4], sp_reg_n_0_[3], sp_reg_n_0_[2]}),
        .S[3:0]({memBAddr[5]_i_3_n_0, memBAddr[5]_i_4_n_0, memBAddr[5]_i_5_n_0, memBAddr[5]_i_6_n_0})
    );
    FDCE memBAddr_reg[6]
    (
        .Q(memBAddr_reg_n_0_[6]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memBAddr[6])
    );
    FDCE memBAddr_reg[7]
    (
        .Q(memBAddr_reg_n_0_[7]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memBAddr[7])
    );
    FDCE memBAddr_reg[8]
    (
        .Q(memBAddr_reg_n_0_[8]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memBAddr[8])
    );
    FDCE memBAddr_reg[9]
    (
        .Q(memBAddr_reg_n_0_[9]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memBAddr[9])
    );
    CARRY4 memBAddr_reg[9]_i_2
    (
        .CI(memBAddr_reg[5]_i_2_n_0),
        .CYINIT(<const0>),
        .CO[3:0]({memBAddr_reg[9]_i_2_n_0, memBAddr_reg[9]_i_2_n_1, memBAddr_reg[9]_i_2_n_2, memBAddr_reg[9]_i_2_n_3}),
        .O[3:0]({memBAddr_reg[9]_i_2_n_4, memBAddr_reg[9]_i_2_n_5, memBAddr_reg[9]_i_2_n_6, memBAddr_reg[9]_i_2_n_7}),
        .DI[3:0]({<const0>, <const0>, <const0>, sp_reg_n_0_[6]}),
        .S[3:0]({memBAddr[9]_i_3_n_0, memBAddr[9]_i_4_n_0, memBAddr[9]_i_5_n_0, memBAddr[9]_i_6_n_0})
    );
    LUT6 memBWriteEnable_i_1
    (
        .O(memBWriteEnable),
        .I0(decodedOpcode_reg_n_0_[4]),
        .I1(decodedOpcode_reg_n_0_[1]),
        .I2(decodedOpcode_reg_n_0_[3]),
        .I3(decodedOpcode_reg_n_0_[2]),
        .I4(decodedOpcode_reg_n_0_[0]),
        .I5(FSM_sequential_state[3]_i_3_n_0)
    );
    FDCE memBWriteEnable_reg
    (
        .Q(memBWriteEnable_reg_n_0),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memBWriteEnable)
    );
    FDCE memBWrite_reg[0]
    (
        .Q(memBWrite[0]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memARead[0])
    );
    FDCE memBWrite_reg[10]
    (
        .Q(memBWrite[10]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memARead[10])
    );
    FDCE memBWrite_reg[11]
    (
        .Q(memBWrite[11]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memARead[11])
    );
    FDCE memBWrite_reg[12]
    (
        .Q(memBWrite[12]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memARead[12])
    );
    FDCE memBWrite_reg[13]
    (
        .Q(memBWrite[13]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memARead[13])
    );
    FDCE memBWrite_reg[14]
    (
        .Q(memBWrite[14]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memARead[14])
    );
    FDCE memBWrite_reg[15]
    (
        .Q(memBWrite[15]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memARead[15])
    );
    FDCE memBWrite_reg[16]
    (
        .Q(memBWrite[16]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memARead[16])
    );
    FDCE memBWrite_reg[17]
    (
        .Q(memBWrite[17]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memARead[17])
    );
    FDCE memBWrite_reg[18]
    (
        .Q(memBWrite[18]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memARead[18])
    );
    FDCE memBWrite_reg[19]
    (
        .Q(memBWrite[19]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memARead[19])
    );
    FDCE memBWrite_reg[1]
    (
        .Q(memBWrite[1]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memARead[1])
    );
    FDCE memBWrite_reg[20]
    (
        .Q(memBWrite[20]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memARead[20])
    );
    FDCE memBWrite_reg[21]
    (
        .Q(memBWrite[21]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memARead[21])
    );
    FDCE memBWrite_reg[22]
    (
        .Q(memBWrite[22]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memARead[22])
    );
    FDCE memBWrite_reg[23]
    (
        .Q(memBWrite[23]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memARead[23])
    );
    FDCE memBWrite_reg[24]
    (
        .Q(memBWrite[24]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memARead[24])
    );
    FDCE memBWrite_reg[25]
    (
        .Q(memBWrite[25]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memARead[25])
    );
    FDCE memBWrite_reg[26]
    (
        .Q(memBWrite[26]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memARead[26])
    );
    FDCE memBWrite_reg[27]
    (
        .Q(memBWrite[27]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memARead[27])
    );
    FDCE memBWrite_reg[28]
    (
        .Q(memBWrite[28]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memARead[28])
    );
    FDCE memBWrite_reg[29]
    (
        .Q(memBWrite[29]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memARead[29])
    );
    FDCE memBWrite_reg[2]
    (
        .Q(memBWrite[2]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memARead[2])
    );
    FDCE memBWrite_reg[30]
    (
        .Q(memBWrite[30]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memARead[30])
    );
    FDCE memBWrite_reg[31]
    (
        .Q(memBWrite[31]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memARead[31])
    );
    FDCE memBWrite_reg[3]
    (
        .Q(memBWrite[3]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memARead[3])
    );
    FDCE memBWrite_reg[4]
    (
        .Q(memBWrite[4]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memARead[4])
    );
    FDCE memBWrite_reg[5]
    (
        .Q(memBWrite[5]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memARead[5])
    );
    FDCE memBWrite_reg[6]
    (
        .Q(memBWrite[6]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memARead[6])
    );
    FDCE memBWrite_reg[7]
    (
        .Q(memBWrite[7]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memARead[7])
    );
    FDCE memBWrite_reg[8]
    (
        .Q(memBWrite[8]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memARead[8])
    );
    FDCE memBWrite_reg[9]
    (
        .Q(memBWrite[9]),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memARead[9])
    );
    IBUF mem_read_IBUF[0]_inst
    (
        .O(mem_read_IBUF[0]),
        .I(mem_read[0])
    );
    IBUF mem_read_IBUF[10]_inst
    (
        .O(mem_read_IBUF[10]),
        .I(mem_read[10])
    );
    IBUF mem_read_IBUF[11]_inst
    (
        .O(mem_read_IBUF[11]),
        .I(mem_read[11])
    );
    IBUF mem_read_IBUF[12]_inst
    (
        .O(mem_read_IBUF[12]),
        .I(mem_read[12])
    );
    IBUF mem_read_IBUF[13]_inst
    (
        .O(mem_read_IBUF[13]),
        .I(mem_read[13])
    );
    IBUF mem_read_IBUF[14]_inst
    (
        .O(mem_read_IBUF[14]),
        .I(mem_read[14])
    );
    IBUF mem_read_IBUF[15]_inst
    (
        .O(mem_read_IBUF[15]),
        .I(mem_read[15])
    );
    IBUF mem_read_IBUF[16]_inst
    (
        .O(mem_read_IBUF[16]),
        .I(mem_read[16])
    );
    IBUF mem_read_IBUF[17]_inst
    (
        .O(mem_read_IBUF[17]),
        .I(mem_read[17])
    );
    IBUF mem_read_IBUF[18]_inst
    (
        .O(mem_read_IBUF[18]),
        .I(mem_read[18])
    );
    IBUF mem_read_IBUF[19]_inst
    (
        .O(mem_read_IBUF[19]),
        .I(mem_read[19])
    );
    IBUF mem_read_IBUF[1]_inst
    (
        .O(mem_read_IBUF[1]),
        .I(mem_read[1])
    );
    IBUF mem_read_IBUF[20]_inst
    (
        .O(mem_read_IBUF[20]),
        .I(mem_read[20])
    );
    IBUF mem_read_IBUF[21]_inst
    (
        .O(mem_read_IBUF[21]),
        .I(mem_read[21])
    );
    IBUF mem_read_IBUF[22]_inst
    (
        .O(mem_read_IBUF[22]),
        .I(mem_read[22])
    );
    IBUF mem_read_IBUF[23]_inst
    (
        .O(mem_read_IBUF[23]),
        .I(mem_read[23])
    );
    IBUF mem_read_IBUF[24]_inst
    (
        .O(mem_read_IBUF[24]),
        .I(mem_read[24])
    );
    IBUF mem_read_IBUF[25]_inst
    (
        .O(mem_read_IBUF[25]),
        .I(mem_read[25])
    );
    IBUF mem_read_IBUF[26]_inst
    (
        .O(mem_read_IBUF[26]),
        .I(mem_read[26])
    );
    IBUF mem_read_IBUF[27]_inst
    (
        .O(mem_read_IBUF[27]),
        .I(mem_read[27])
    );
    IBUF mem_read_IBUF[28]_inst
    (
        .O(mem_read_IBUF[28]),
        .I(mem_read[28])
    );
    IBUF mem_read_IBUF[29]_inst
    (
        .O(mem_read_IBUF[29]),
        .I(mem_read[29])
    );
    IBUF mem_read_IBUF[2]_inst
    (
        .O(mem_read_IBUF[2]),
        .I(mem_read[2])
    );
    IBUF mem_read_IBUF[30]_inst
    (
        .O(mem_read_IBUF[30]),
        .I(mem_read[30])
    );
    IBUF mem_read_IBUF[31]_inst
    (
        .O(mem_read_IBUF[31]),
        .I(mem_read[31])
    );
    IBUF mem_read_IBUF[3]_inst
    (
        .O(mem_read_IBUF[3]),
        .I(mem_read[3])
    );
    IBUF mem_read_IBUF[4]_inst
    (
        .O(mem_read_IBUF[4]),
        .I(mem_read[4])
    );
    IBUF mem_read_IBUF[5]_inst
    (
        .O(mem_read_IBUF[5]),
        .I(mem_read[5])
    );
    IBUF mem_read_IBUF[6]_inst
    (
        .O(mem_read_IBUF[6]),
        .I(mem_read[6])
    );
    IBUF mem_read_IBUF[7]_inst
    (
        .O(mem_read_IBUF[7]),
        .I(mem_read[7])
    );
    IBUF mem_read_IBUF[8]_inst
    (
        .O(mem_read_IBUF[8]),
        .I(mem_read[8])
    );
    IBUF mem_read_IBUF[9]_inst
    (
        .O(mem_read_IBUF[9]),
        .I(mem_read[9])
    );
    OBUF mem_writeMask_OBUF[0]_inst
    (
        .O(mem_writeMask[0]),
        .I(<const1>)
    );
    OBUF mem_writeMask_OBUF[1]_inst
    (
        .O(mem_writeMask[1]),
        .I(<const1>)
    );
    OBUF mem_writeMask_OBUF[2]_inst
    (
        .O(mem_writeMask[2]),
        .I(<const1>)
    );
    OBUF mem_writeMask_OBUF[3]_inst
    (
        .O(mem_writeMask[3]),
        .I(<const1>)
    );
    LUT1 mem_write[31]_i_1
    (
        .O(mem_write[31]_i_1_n_0),
        .I0(areset_IBUF)
    );
    OBUF mem_write_OBUF[0]_inst
    (
        .O(mem_write[0]),
        .I(mem_write_OBUF[0])
    );
    OBUF mem_write_OBUF[10]_inst
    (
        .O(mem_write[10]),
        .I(mem_write_OBUF[10])
    );
    OBUF mem_write_OBUF[11]_inst
    (
        .O(mem_write[11]),
        .I(mem_write_OBUF[11])
    );
    OBUF mem_write_OBUF[12]_inst
    (
        .O(mem_write[12]),
        .I(mem_write_OBUF[12])
    );
    OBUF mem_write_OBUF[13]_inst
    (
        .O(mem_write[13]),
        .I(mem_write_OBUF[13])
    );
    OBUF mem_write_OBUF[14]_inst
    (
        .O(mem_write[14]),
        .I(mem_write_OBUF[14])
    );
    OBUF mem_write_OBUF[15]_inst
    (
        .O(mem_write[15]),
        .I(mem_write_OBUF[15])
    );
    OBUF mem_write_OBUF[16]_inst
    (
        .O(mem_write[16]),
        .I(mem_write_OBUF[16])
    );
    OBUF mem_write_OBUF[17]_inst
    (
        .O(mem_write[17]),
        .I(mem_write_OBUF[17])
    );
    OBUF mem_write_OBUF[18]_inst
    (
        .O(mem_write[18]),
        .I(mem_write_OBUF[18])
    );
    OBUF mem_write_OBUF[19]_inst
    (
        .O(mem_write[19]),
        .I(mem_write_OBUF[19])
    );
    OBUF mem_write_OBUF[1]_inst
    (
        .O(mem_write[1]),
        .I(mem_write_OBUF[1])
    );
    OBUF mem_write_OBUF[20]_inst
    (
        .O(mem_write[20]),
        .I(mem_write_OBUF[20])
    );
    OBUF mem_write_OBUF[21]_inst
    (
        .O(mem_write[21]),
        .I(mem_write_OBUF[21])
    );
    OBUF mem_write_OBUF[22]_inst
    (
        .O(mem_write[22]),
        .I(mem_write_OBUF[22])
    );
    OBUF mem_write_OBUF[23]_inst
    (
        .O(mem_write[23]),
        .I(mem_write_OBUF[23])
    );
    OBUF mem_write_OBUF[24]_inst
    (
        .O(mem_write[24]),
        .I(mem_write_OBUF[24])
    );
    OBUF mem_write_OBUF[25]_inst
    (
        .O(mem_write[25]),
        .I(mem_write_OBUF[25])
    );
    OBUF mem_write_OBUF[26]_inst
    (
        .O(mem_write[26]),
        .I(mem_write_OBUF[26])
    );
    OBUF mem_write_OBUF[27]_inst
    (
        .O(mem_write[27]),
        .I(mem_write_OBUF[27])
    );
    OBUF mem_write_OBUF[28]_inst
    (
        .O(mem_write[28]),
        .I(mem_write_OBUF[28])
    );
    OBUF mem_write_OBUF[29]_inst
    (
        .O(mem_write[29]),
        .I(mem_write_OBUF[29])
    );
    OBUF mem_write_OBUF[2]_inst
    (
        .O(mem_write[2]),
        .I(mem_write_OBUF[2])
    );
    OBUF mem_write_OBUF[30]_inst
    (
        .O(mem_write[30]),
        .I(mem_write_OBUF[30])
    );
    OBUF mem_write_OBUF[31]_inst
    (
        .O(mem_write[31]),
        .I(mem_write_OBUF[31])
    );
    OBUF mem_write_OBUF[3]_inst
    (
        .O(mem_write[3]),
        .I(mem_write_OBUF[3])
    );
    OBUF mem_write_OBUF[4]_inst
    (
        .O(mem_write[4]),
        .I(mem_write_OBUF[4])
    );
    OBUF mem_write_OBUF[5]_inst
    (
        .O(mem_write[5]),
        .I(mem_write_OBUF[5])
    );
    OBUF mem_write_OBUF[6]_inst
    (
        .O(mem_write[6]),
        .I(mem_write_OBUF[6])
    );
    OBUF mem_write_OBUF[7]_inst
    (
        .O(mem_write[7]),
        .I(mem_write_OBUF[7])
    );
    OBUF mem_write_OBUF[8]_inst
    (
        .O(mem_write[8]),
        .I(mem_write_OBUF[8])
    );
    OBUF mem_write_OBUF[9]_inst
    (
        .O(mem_write[9]),
        .I(mem_write_OBUF[9])
    );
    FDRE mem_write_reg[0]
    (
        .Q(mem_write_OBUF[0]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memBRead[0]),
        .R(<const0>)
    );
    FDRE mem_write_reg[10]
    (
        .Q(mem_write_OBUF[10]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memBRead[10]),
        .R(<const0>)
    );
    FDRE mem_write_reg[11]
    (
        .Q(mem_write_OBUF[11]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memBRead[11]),
        .R(<const0>)
    );
    FDRE mem_write_reg[12]
    (
        .Q(mem_write_OBUF[12]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memBRead[12]),
        .R(<const0>)
    );
    FDRE mem_write_reg[13]
    (
        .Q(mem_write_OBUF[13]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memBRead[13]),
        .R(<const0>)
    );
    FDRE mem_write_reg[14]
    (
        .Q(mem_write_OBUF[14]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memBRead[14]),
        .R(<const0>)
    );
    FDRE mem_write_reg[15]
    (
        .Q(mem_write_OBUF[15]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memBRead[15]),
        .R(<const0>)
    );
    FDRE mem_write_reg[16]
    (
        .Q(mem_write_OBUF[16]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memBRead[16]),
        .R(<const0>)
    );
    FDRE mem_write_reg[17]
    (
        .Q(mem_write_OBUF[17]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memBRead[17]),
        .R(<const0>)
    );
    FDRE mem_write_reg[18]
    (
        .Q(mem_write_OBUF[18]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memBRead[18]),
        .R(<const0>)
    );
    FDRE mem_write_reg[19]
    (
        .Q(mem_write_OBUF[19]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memBRead[19]),
        .R(<const0>)
    );
    FDRE mem_write_reg[1]
    (
        .Q(mem_write_OBUF[1]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memBRead[1]),
        .R(<const0>)
    );
    FDRE mem_write_reg[20]
    (
        .Q(mem_write_OBUF[20]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memBRead[20]),
        .R(<const0>)
    );
    FDRE mem_write_reg[21]
    (
        .Q(mem_write_OBUF[21]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memBRead[21]),
        .R(<const0>)
    );
    FDRE mem_write_reg[22]
    (
        .Q(mem_write_OBUF[22]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memBRead[22]),
        .R(<const0>)
    );
    FDRE mem_write_reg[23]
    (
        .Q(mem_write_OBUF[23]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memBRead[23]),
        .R(<const0>)
    );
    FDRE mem_write_reg[24]
    (
        .Q(mem_write_OBUF[24]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memBRead[24]),
        .R(<const0>)
    );
    FDRE mem_write_reg[25]
    (
        .Q(mem_write_OBUF[25]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memBRead[25]),
        .R(<const0>)
    );
    FDRE mem_write_reg[26]
    (
        .Q(mem_write_OBUF[26]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memBRead[26]),
        .R(<const0>)
    );
    FDRE mem_write_reg[27]
    (
        .Q(mem_write_OBUF[27]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memBRead[27]),
        .R(<const0>)
    );
    FDRE mem_write_reg[28]
    (
        .Q(mem_write_OBUF[28]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memBRead[28]),
        .R(<const0>)
    );
    FDRE mem_write_reg[29]
    (
        .Q(mem_write_OBUF[29]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memBRead[29]),
        .R(<const0>)
    );
    FDRE mem_write_reg[2]
    (
        .Q(mem_write_OBUF[2]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memBRead[2]),
        .R(<const0>)
    );
    FDRE mem_write_reg[30]
    (
        .Q(mem_write_OBUF[30]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memBRead[30]),
        .R(<const0>)
    );
    FDRE mem_write_reg[31]
    (
        .Q(mem_write_OBUF[31]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memBRead[31]),
        .R(<const0>)
    );
    FDRE mem_write_reg[3]
    (
        .Q(mem_write_OBUF[3]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memBRead[3]),
        .R(<const0>)
    );
    FDRE mem_write_reg[4]
    (
        .Q(mem_write_OBUF[4]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memBRead[4]),
        .R(<const0>)
    );
    FDRE mem_write_reg[5]
    (
        .Q(mem_write_OBUF[5]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memBRead[5]),
        .R(<const0>)
    );
    FDRE mem_write_reg[6]
    (
        .Q(mem_write_OBUF[6]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memBRead[6]),
        .R(<const0>)
    );
    FDRE mem_write_reg[7]
    (
        .Q(mem_write_OBUF[7]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memBRead[7]),
        .R(<const0>)
    );
    FDRE mem_write_reg[8]
    (
        .Q(mem_write_OBUF[8]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memBRead[8]),
        .R(<const0>)
    );
    FDRE mem_write_reg[9]
    (
        .Q(mem_write_OBUF[9]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memBRead[9]),
        .R(<const0>)
    );
    dualport_ram memory
    (
        .FSM_sequential_state_reg[0](FSM_sequential_state[2]_i_3_n_0),
        .FSM_sequential_state_reg[1](FSM_sequential_state[3]_i_5_n_0),
        .FSM_sequential_state_reg[1]_0(decodedOpcode[4]_i_2_n_0),
        .FSM_sequential_state_reg[2](FSM_sequential_state[1]_i_3_n_0),
        .FSM_sequential_state_reg[3](FSM_sequential_state[3]_i_3_n_0),
        .clk_IBUF_BUFG(clk_IBUF_BUFG),
        .decodedOpcode_reg[0](pc[9]_i_2_n_0),
        .decodedOpcode_reg[0]_0(pc[9]_i_3_n_0),
        .decodedOpcode_reg[0]_1(pc[9]_i_4_n_0),
        .decodedOpcode_reg[0]_2(pc[14]_i_5_n_0),
        .decodedOpcode_reg[0]_3(memAAddr[2]_i_3_n_0),
        .decodedOpcode_reg[0]_4(sp[14]_i_8_n_0),
        .decodedOpcode_reg[1](memAAddr[14]_i_5_n_0),
        .decodedOpcode_reg[2](out_mem_readEnable_i_2_n_0),
        .decodedOpcode_reg[2]_0(memAWrite[31]_i_4_n_0),
        .decodedOpcode_reg[2]_1(sp[14]_i_4_n_0),
        .decodedOpcode_reg[2]_10(memAAddr[7]_i_4_n_0),
        .decodedOpcode_reg[2]_11(memAAddr[8]_i_4_n_0),
        .decodedOpcode_reg[2]_12(memAAddr[9]_i_4_n_0),
        .decodedOpcode_reg[2]_13(memAAddr[10]_i_4_n_0),
        .decodedOpcode_reg[2]_14(memAAddr[11]_i_4_n_0),
        .decodedOpcode_reg[2]_15(memAAddr[12]_i_4_n_0),
        .decodedOpcode_reg[2]_16(memAAddr[13]_i_4_n_0),
        .decodedOpcode_reg[2]_17(memAAddr[14]_i_6_n_0),
        .decodedOpcode_reg[2]_2(sp[14]_i_6_n_0),
        .decodedOpcode_reg[2]_3(pc[5]_i_3_n_0),
        .decodedOpcode_reg[2]_4(pc[14]_i_3_n_0),
        .decodedOpcode_reg[2]_5(memAAddr[2]_i_4_n_0),
        .decodedOpcode_reg[2]_6(memAAddr[3]_i_4_n_0),
        .decodedOpcode_reg[2]_7(memAAddr[4]_i_4_n_0),
        .decodedOpcode_reg[2]_8(memAAddr[5]_i_4_n_0),
        .decodedOpcode_reg[2]_9(memAAddr[6]_i_4_n_0),
        .decodedOpcode_reg[3](memAWrite[14]_i_7_n_0),
        .decodedOpcode_reg[3]_0(memAWrite[13]_i_7_n_0),
        .decodedOpcode_reg[3]_1(memAWrite[12]_i_7_n_0),
        .decodedOpcode_reg[3]_10(memAWrite[3]_i_5_n_0),
        .decodedOpcode_reg[3]_11(memAWrite[2]_i_5_n_0),
        .decodedOpcode_reg[3]_12(pc[5]_i_4_n_0),
        .decodedOpcode_reg[3]_2(memAWrite[11]_i_7_n_0),
        .decodedOpcode_reg[3]_3(memAWrite[10]_i_7_n_0),
        .decodedOpcode_reg[3]_4(memAWrite[9]_i_7_n_0),
        .decodedOpcode_reg[3]_5(memAWrite[8]_i_7_n_0),
        .decodedOpcode_reg[3]_6(memAWrite[7]_i_7_n_0),
        .decodedOpcode_reg[3]_7(memAWrite[6]_i_5_n_0),
        .decodedOpcode_reg[3]_8(memAWrite[5]_i_5_n_0),
        .decodedOpcode_reg[3]_9(memAWrite[4]_i_5_n_0),
        .decodedOpcode_reg[4]_0(sp[2]_i_2_n_0),
        .decodedOpcode_reg[4]_1(memAAddr[14]_i_4_n_0),
        .idim_flag(idim_flag),
        .inInterrupt_reg(decodedOpcode[4]_i_5_n_0),
        .in_mem_busy_IBUF(in_mem_busy_IBUF),
        .memAWriteEnable(memAWriteEnable_reg_n_0),
        .memBWriteEnable(memBWriteEnable_reg_n_0),
        .opcode_reg[0](memory_n_148),
        .opcode_reg[0]_0(memAWrite[0]_i_4_n_0),
        .opcode_reg[0]_1(pc[5]_i_2_n_0),
        .opcode_reg[1](memory_n_149),
        .opcode_reg[1]_0(memAWrite[1]_i_4_n_0),
        .opcode_reg[2](memory_n_150),
        .opcode_reg[3](memory_n_151),
        .opcode_reg[4](memory_n_152),
        .opcode_reg[5](memory_n_42),
        .opcode_reg[6](memory_n_41),
        .out_mem_readEnable_reg(memory_n_3),
        .pc_reg[10](memAWrite[10]_i_4_n_0),
        .pc_reg[11](memAWrite[11]_i_4_n_0),
        .pc_reg[12](memAWrite[12]_i_4_n_0),
        .pc_reg[13](memAWrite[13]_i_4_n_0),
        .pc_reg[14]_0(memAWrite[14]_i_4_n_0),
        .pc_reg[2](memAWrite[2]_i_4_n_0),
        .pc_reg[3](memAWrite[3]_i_4_n_0),
        .pc_reg[4](memAWrite[4]_i_4_n_0),
        .pc_reg[5](memAWrite[5]_i_4_n_0),
        .pc_reg[6](memAWrite[6]_i_4_n_0),
        .pc_reg[7](memAWrite[7]_i_4_n_0),
        .pc_reg[8](memAWrite[8]_i_4_n_0),
        .pc_reg[9](memAWrite[9]_i_4_n_0),
        .D[2:0]({memory_n_0, memory_n_1, memory_n_2}),
        .O[3:0]({sp_reg[14]_i_7_n_4, sp_reg[14]_i_7_n_5, sp_reg[14]_i_7_n_6, sp_reg[14]_i_7_n_7}),
        .Q[4:0]({decodedOpcode_reg_n_0_[4], decodedOpcode_reg_n_0_[3], decodedOpcode_reg_n_0_[2], decodedOpcode_reg_n_0_[1], decodedOpcode_reg_n_0_[0]}),
        .data2[11:0]({sp_reg[14]_i_5_n_4, sp_reg[14]_i_5_n_5, sp_reg[14]_i_5_n_6, sp_reg[14]_i_5_n_7, sp_reg[10]_i_3_n_4, sp_reg[10]_i_3_n_5, sp_reg[10]_i_3_n_6, sp_reg[10]_i_3_n_7, sp_reg[6]_i_3_n_4, sp_reg[6]_i_3_n_5, sp_reg[6]_i_3_n_6, sp_reg[6]_i_3_n_7}),
        .decodedOpcode_reg[4][4:0]({decodedOpcode[4], decodedOpcode[3], decodedOpcode[2], decodedOpcode[1], decodedOpcode[0]}),
        .memAAddr_reg[14][12:0]({memAAddr[14], memAAddr[13], memAAddr[12], memAAddr[11], memAAddr[10], memAAddr[9], memAAddr[8], memAAddr[7], memAAddr[6], memAAddr[5], memAAddr[4], memAAddr[3], memAAddr[2]}),
        .memAAddr_reg[14]_0[12:0]({memAAddr_reg_n_0_[14], memAAddr_reg_n_0_[13], memAAddr_reg_n_0_[12], memAAddr_reg_n_0_[11], memAAddr_reg_n_0_[10], memAAddr_reg_n_0_[9], memAAddr_reg_n_0_[8], memAAddr_reg_n_0_[7], memAAddr_reg_n_0_[6], memAAddr_reg_n_0_[5], memAAddr_reg_n_0_[4], memAAddr_reg_n_0_[3], memAAddr_reg_n_0_[2]}),
        .memARead[31:0]({memARead[31], memARead[30], memARead[29], memARead[28], memARead[27], memARead[26], memARead[25], memARead[24], memARead[23], memARead[22], memARead[21], memARead[20], memARead[19], memARead[18], memARead[17], memARead[16], memARead[15], memARead[14], memARead[13], memARead[12], memARead[11], memARead[10], memARead[9], memARead[8], memARead[7], memARead[6], memARead[5], memARead[4], memARead[3], memARead[2], memARead[1], memARead[0]}),
        .memAWrite_reg[31][31:0]({memAWrite[31], memAWrite[30], memAWrite[29], memAWrite[28], memAWrite[27], memAWrite[26], memAWrite[25], memAWrite[24], memAWrite[23], memAWrite[22], memAWrite[21], memAWrite[20], memAWrite[19], memAWrite[18], memAWrite[17], memAWrite[16], memAWrite[15], memAWrite[14], memAWrite[13], memAWrite[12], memAWrite[11], memAWrite[10], memAWrite[9], memAWrite[8], memAWrite[7], memAWrite[6], memAWrite[5], memAWrite[4], memAWrite[3], memAWrite[2], memAWrite[1], memAWrite[0]}),
        .memAWrite_reg[31]_0[31:0]({memAWrite_reg_n_0_[31], memAWrite_reg_n_0_[30], memAWrite_reg_n_0_[29], memAWrite_reg_n_0_[28], memAWrite_reg_n_0_[27], memAWrite_reg_n_0_[26], memAWrite_reg_n_0_[25], memAWrite_reg_n_0_[24], memAWrite_reg_n_0_[23], memAWrite_reg_n_0_[22], memAWrite_reg_n_0_[21], memAWrite_reg_n_0_[20], memAWrite_reg_n_0_[19], memAWrite_reg_n_0_[18], memAWrite_reg_n_0_[17], memAWrite_reg_n_0_[16], memAWrite_reg_n_0_[15], memAWrite_reg_n_0_[14], memAWrite_reg_n_0_[13], memAWrite_reg_n_0_[12], memAWrite_reg_n_0_[11], memAWrite_reg_n_0_[10], memAWrite_reg_n_0_[9], memAWrite_reg_n_0_[8], memAWrite_reg_n_0_[7], memAWrite_reg_n_0_[6], memAWrite_reg_n_0_[5], memAWrite_reg_n_0_[4], memAWrite_reg_n_0_[3], memAWrite_reg_n_0_[2], memAWrite_reg_n_0_[1], memAWrite_reg_n_0_[0]}),
        .memBAddr_reg[14][12:0]({memBAddr_reg_n_0_[14], memBAddr_reg_n_0_[13], memBAddr_reg_n_0_[12], memBAddr_reg_n_0_[11], memBAddr_reg_n_0_[10], memBAddr_reg_n_0_[9], memBAddr_reg_n_0_[8], memBAddr_reg_n_0_[7], memBAddr_reg_n_0_[6], memBAddr_reg_n_0_[5], memBAddr_reg_n_0_[4], memBAddr_reg_n_0_[3], memBAddr_reg_n_0_[2]}),
        .memBRead[31:0]({memBRead[31], memBRead[30], memBRead[29], memBRead[28], memBRead[27], memBRead[26], memBRead[25], memBRead[24], memBRead[23], memBRead[22], memBRead[21], memBRead[20], memBRead[19], memBRead[18], memBRead[17], memBRead[16], memBRead[15], memBRead[14], memBRead[13], memBRead[12], memBRead[11], memBRead[10], memBRead[9], memBRead[8], memBRead[7], memBRead[6], memBRead[5], memBRead[4], memBRead[3], memBRead[2], memBRead[1], memBRead[0]}),
        .memBWrite_reg[31][31:0]({memBWrite[31], memBWrite[30], memBWrite[29], memBWrite[28], memBWrite[27], memBWrite[26], memBWrite[25], memBWrite[24], memBWrite[23], memBWrite[22], memBWrite[21], memBWrite[20], memBWrite[19], memBWrite[18], memBWrite[17], memBWrite[16], memBWrite[15], memBWrite[14], memBWrite[13], memBWrite[12], memBWrite[11], memBWrite[10], memBWrite[9], memBWrite[8], memBWrite[7], memBWrite[6], memBWrite[5], memBWrite[4], memBWrite[3], memBWrite[2], memBWrite[1], memBWrite[0]}),
        .mem_read_IBUF[31:0]({mem_read_IBUF[31], mem_read_IBUF[30], mem_read_IBUF[29], mem_read_IBUF[28], mem_read_IBUF[27], mem_read_IBUF[26], mem_read_IBUF[25], mem_read_IBUF[24], mem_read_IBUF[23], mem_read_IBUF[22], mem_read_IBUF[21], mem_read_IBUF[20], mem_read_IBUF[19], mem_read_IBUF[18], mem_read_IBUF[17], mem_read_IBUF[16], mem_read_IBUF[15], mem_read_IBUF[14], mem_read_IBUF[13], mem_read_IBUF[12], mem_read_IBUF[11], mem_read_IBUF[10], mem_read_IBUF[9], mem_read_IBUF[8], mem_read_IBUF[7], mem_read_IBUF[6], mem_read_IBUF[5], mem_read_IBUF[4], mem_read_IBUF[3], mem_read_IBUF[2], mem_read_IBUF[1], mem_read_IBUF[0]}),
        .opcode_reg[6]_0[4:0]({opcode_reg_n_0_[6], opcode_reg_n_0_[4], opcode_reg_n_0_[3], opcode_reg_n_0_[2], opcode_reg_n_0_[1]}),
        .out[3:0]({FSM_sequential_state_reg_n_0_[3], FSM_sequential_state_reg_n_0_[2], FSM_sequential_state_reg_n_0_[1], FSM_sequential_state_reg_n_0_[0]}),
        .pc_reg[14][14:0]({pc[14], pc[13], pc[12], pc[11], pc[10], pc[9], pc[8], pc[7], pc[6], pc[5], pc[4], pc[3], pc[2], pc[1], pc[0]}),
        .pc_reg[14]_1[13:0]({data2[14], data2[13], data2[12], data2[11], data2[10], data2[9], data2[8], data2[7], data2[6], data2[5], data2[4], data2[3], data2[2], data2[1]}),
        .pc_reg[1][1:0]({data0[1], data0[0]}),
        .sp_reg[10][3:0]({sp_reg[10]_i_4_n_4, sp_reg[10]_i_4_n_5, sp_reg[10]_i_4_n_6, sp_reg[10]_i_4_n_7}),
        .sp_reg[14][12:0]({sp[14], sp[13], sp[12], sp[11], sp[10], sp[9], sp[8], sp[7], sp[6], sp[5], sp[4], sp[3], sp[2]}),
        .sp_reg[14]_0[12:0]({sp_reg_n_0_[14], sp_reg_n_0_[13], sp_reg_n_0_[12], sp_reg_n_0_[11], sp_reg_n_0_[10], sp_reg_n_0_[9], sp_reg_n_0_[8], sp_reg_n_0_[7], sp_reg_n_0_[6], sp_reg_n_0_[5], sp_reg_n_0_[4], sp_reg_n_0_[3], sp_reg_n_0_[2]}),
        .sp_reg[2][3:0]({sp_reg[6]_i_4_n_4, sp_reg[6]_i_4_n_5, sp_reg[6]_i_4_n_6, sp_reg[6]_i_4_n_7})
    );
    FDRE opcode_reg[0]
    (
        .Q(opcode_reg_n_0_[0]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memory_n_148),
        .R(<const0>)
    );
    FDRE opcode_reg[1]
    (
        .Q(opcode_reg_n_0_[1]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memory_n_149),
        .R(<const0>)
    );
    FDRE opcode_reg[2]
    (
        .Q(opcode_reg_n_0_[2]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memory_n_150),
        .R(<const0>)
    );
    FDRE opcode_reg[3]
    (
        .Q(opcode_reg_n_0_[3]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memory_n_151),
        .R(<const0>)
    );
    FDRE opcode_reg[4]
    (
        .Q(opcode_reg_n_0_[4]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memory_n_152),
        .R(<const0>)
    );
    FDRE opcode_reg[5]
    (
        .Q(opcode_reg_n_0_[5]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memory_n_42),
        .R(<const0>)
    );
    FDRE opcode_reg[6]
    (
        .Q(opcode_reg_n_0_[6]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memory_n_41),
        .R(<const0>)
    );
    OBUF out_mem_addr_OBUF[0]_inst
    (
        .O(out_mem_addr[0]),
        .I(out_mem_addr_OBUF[0])
    );
    OBUF out_mem_addr_OBUF[10]_inst
    (
        .O(out_mem_addr[10]),
        .I(out_mem_addr_OBUF[10])
    );
    OBUF out_mem_addr_OBUF[11]_inst
    (
        .O(out_mem_addr[11]),
        .I(out_mem_addr_OBUF[11])
    );
    OBUF out_mem_addr_OBUF[12]_inst
    (
        .O(out_mem_addr[12]),
        .I(out_mem_addr_OBUF[12])
    );
    OBUF out_mem_addr_OBUF[13]_inst
    (
        .O(out_mem_addr[13]),
        .I(out_mem_addr_OBUF[13])
    );
    OBUF out_mem_addr_OBUF[14]_inst
    (
        .O(out_mem_addr[14]),
        .I(out_mem_addr_OBUF[14])
    );
    OBUF out_mem_addr_OBUF[15]_inst
    (
        .O(out_mem_addr[15]),
        .I(out_mem_addr_OBUF[15])
    );
    OBUF out_mem_addr_OBUF[1]_inst
    (
        .O(out_mem_addr[1]),
        .I(out_mem_addr_OBUF[1])
    );
    OBUF out_mem_addr_OBUF[2]_inst
    (
        .O(out_mem_addr[2]),
        .I(out_mem_addr_OBUF[2])
    );
    OBUF out_mem_addr_OBUF[3]_inst
    (
        .O(out_mem_addr[3]),
        .I(out_mem_addr_OBUF[3])
    );
    OBUF out_mem_addr_OBUF[4]_inst
    (
        .O(out_mem_addr[4]),
        .I(out_mem_addr_OBUF[4])
    );
    OBUF out_mem_addr_OBUF[5]_inst
    (
        .O(out_mem_addr[5]),
        .I(out_mem_addr_OBUF[5])
    );
    OBUF out_mem_addr_OBUF[6]_inst
    (
        .O(out_mem_addr[6]),
        .I(out_mem_addr_OBUF[6])
    );
    OBUF out_mem_addr_OBUF[7]_inst
    (
        .O(out_mem_addr[7]),
        .I(out_mem_addr_OBUF[7])
    );
    OBUF out_mem_addr_OBUF[8]_inst
    (
        .O(out_mem_addr[8]),
        .I(out_mem_addr_OBUF[8])
    );
    OBUF out_mem_addr_OBUF[9]_inst
    (
        .O(out_mem_addr[9]),
        .I(out_mem_addr_OBUF[9])
    );
    FDRE out_mem_addr_reg[0]
    (
        .Q(out_mem_addr_OBUF[0]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memARead[0]),
        .R(<const0>)
    );
    FDRE out_mem_addr_reg[10]
    (
        .Q(out_mem_addr_OBUF[10]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memARead[10]),
        .R(<const0>)
    );
    FDRE out_mem_addr_reg[11]
    (
        .Q(out_mem_addr_OBUF[11]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memARead[11]),
        .R(<const0>)
    );
    FDRE out_mem_addr_reg[12]
    (
        .Q(out_mem_addr_OBUF[12]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memARead[12]),
        .R(<const0>)
    );
    FDRE out_mem_addr_reg[13]
    (
        .Q(out_mem_addr_OBUF[13]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memARead[13]),
        .R(<const0>)
    );
    FDRE out_mem_addr_reg[14]
    (
        .Q(out_mem_addr_OBUF[14]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memARead[14]),
        .R(<const0>)
    );
    FDRE out_mem_addr_reg[15]
    (
        .Q(out_mem_addr_OBUF[15]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memARead[15]),
        .R(<const0>)
    );
    FDRE out_mem_addr_reg[1]
    (
        .Q(out_mem_addr_OBUF[1]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memARead[1]),
        .R(<const0>)
    );
    FDRE out_mem_addr_reg[2]
    (
        .Q(out_mem_addr_OBUF[2]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memARead[2]),
        .R(<const0>)
    );
    FDRE out_mem_addr_reg[3]
    (
        .Q(out_mem_addr_OBUF[3]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memARead[3]),
        .R(<const0>)
    );
    FDRE out_mem_addr_reg[4]
    (
        .Q(out_mem_addr_OBUF[4]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memARead[4]),
        .R(<const0>)
    );
    FDRE out_mem_addr_reg[5]
    (
        .Q(out_mem_addr_OBUF[5]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memARead[5]),
        .R(<const0>)
    );
    FDRE out_mem_addr_reg[6]
    (
        .Q(out_mem_addr_OBUF[6]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memARead[6]),
        .R(<const0>)
    );
    FDRE out_mem_addr_reg[7]
    (
        .Q(out_mem_addr_OBUF[7]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memARead[7]),
        .R(<const0>)
    );
    FDRE out_mem_addr_reg[8]
    (
        .Q(out_mem_addr_OBUF[8]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memARead[8]),
        .R(<const0>)
    );
    FDRE out_mem_addr_reg[9]
    (
        .Q(out_mem_addr_OBUF[9]),
        .C(clk_IBUF_BUFG),
        .CE(mem_write[31]_i_1_n_0),
        .D(memARead[9]),
        .R(<const0>)
    );
    OBUF out_mem_readEnable_OBUF_inst
    (
        .O(out_mem_readEnable),
        .I(out_mem_readEnable_OBUF)
    );
    LUT3 out_mem_readEnable_i_2
    (
        .O(out_mem_readEnable_i_2_n_0),
        .I0(decodedOpcode_reg_n_0_[2]),
        .I1(decodedOpcode_reg_n_0_[3]),
        .I2(decodedOpcode_reg_n_0_[0])
    );
    FDCE out_mem_readEnable_reg
    (
        .Q(out_mem_readEnable_OBUF),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(memory_n_3)
    );
    OBUF out_mem_writeEnable_OBUF_inst
    (
        .O(out_mem_writeEnable),
        .I(out_mem_writeEnable_OBUF)
    );
    LUT4 out_mem_writeEnable_i_1
    (
        .O(out_mem_writeEnable_i_1_n_0),
        .I0(FSM_sequential_state_reg_n_0_[3]),
        .I1(FSM_sequential_state_reg_n_0_[0]),
        .I2(FSM_sequential_state_reg_n_0_[1]),
        .I3(FSM_sequential_state_reg_n_0_[2])
    );
    FDCE out_mem_writeEnable_reg
    (
        .Q(out_mem_writeEnable_OBUF),
        .C(clk_IBUF_BUFG),
        .CE(<const1>),
        .CLR(areset_IBUF),
        .D(out_mem_writeEnable_i_1_n_0)
    );
    LUT1 pc[12]_i_3
    (
        .O(pc[12]_i_3_n_0),
        .I0(p_1_in[10])
    );
    LUT1 pc[12]_i_4
    (
        .O(pc[12]_i_4_n_0),
        .I0(p_1_in[9])
    );
    LUT1 pc[12]_i_5
    (
        .O(pc[12]_i_5_n_0),
        .I0(p_1_in[8])
    );
    LUT1 pc[12]_i_6
    (
        .O(pc[12]_i_6_n_0),
        .I0(p_1_in[7])
    );
    LUT4 pc[14]_i_1
    (
        .O(pc[14]_i_1_n_0),
        .I0(FSM_sequential_state_reg_n_0_[1]),
        .I1(FSM_sequential_state_reg_n_0_[2]),
        .I2(FSM_sequential_state_reg_n_0_[0]),
        .I3(FSM_sequential_state_reg_n_0_[3])
    );
    LUT5 pc[14]_i_3
    (
        .O(pc[14]_i_3_n_0),
        .I0(decodedOpcode_reg_n_0_[2]),
        .I1(decodedOpcode_reg_n_0_[0]),
        .I2(decodedOpcode_reg_n_0_[4]),
        .I3(decodedOpcode_reg_n_0_[1]),
        .I4(decodedOpcode_reg_n_0_[3])
    );
    LUT5 pc[14]_i_5
    (
        .O(pc[14]_i_5_n_0),
        .I0(decodedOpcode_reg_n_0_[0]),
        .I1(decodedOpcode_reg_n_0_[1]),
        .I2(decodedOpcode_reg_n_0_[4]),
        .I3(decodedOpcode_reg_n_0_[3]),
        .I4(decodedOpcode_reg_n_0_[2])
    );
    LUT1 pc[14]_i_6
    (
        .O(pc[14]_i_6_n_0),
        .I0(p_1_in[12])
    );
    LUT1 pc[14]_i_7
    (
        .O(pc[14]_i_7_n_0),
        .I0(p_1_in[11])
    );
    LUT1 pc[4]_i_3
    (
        .O(pc[4]_i_3_n_0),
        .I0(p_1_in[2])
    );
    LUT1 pc[4]_i_4
    (
        .O(pc[4]_i_4_n_0),
        .I0(p_1_in[1])
    );
    LUT1 pc[4]_i_5
    (
        .O(pc[4]_i_5_n_0),
        .I0(p_1_in[0])
    );
    LUT1 pc[4]_i_6
    (
        .O(pc[4]_i_6_n_0),
        .I0(data0[1])
    );
    LUT6 pc[5]_i_2
    (
        .O(pc[5]_i_2_n_0),
        .I0(pc[5]_i_5_n_0),
        .I1(opcode_reg_n_0_[0]),
        .I2(decodedOpcode_reg_n_0_[3]),
        .I3(decodedOpcode_reg_n_0_[2]),
        .I4(decodedOpcode_reg_n_0_[0]),
        .I5(data2[5])
    );
    LUT6 pc[5]_i_3
    (
        .O(pc[5]_i_3_n_0),
        .I0(decodedOpcode_reg_n_0_[2]),
        .I1(decodedOpcode_reg_n_0_[1]),
        .I2(decodedOpcode_reg_n_0_[4]),
        .I3(decodedOpcode_reg_n_0_[3]),
        .I4(data2[5]),
        .I5(decodedOpcode_reg_n_0_[0])
    );
    LUT4 pc[5]_i_4
    (
        .O(pc[5]_i_4_n_0),
        .I0(decodedOpcode_reg_n_0_[3]),
        .I1(decodedOpcode_reg_n_0_[2]),
        .I2(decodedOpcode_reg_n_0_[1]),
        .I3(decodedOpcode_reg_n_0_[4])
    );
    LUT2 pc[5]_i_5
    (
        .O(pc[5]_i_5_n_0),
        .I0(decodedOpcode_reg_n_0_[4]),
        .I1(decodedOpcode_reg_n_0_[1])
    );
    LUT1 pc[8]_i_3
    (
        .O(pc[8]_i_3_n_0),
        .I0(p_1_in[6])
    );
    LUT1 pc[8]_i_4
    (
        .O(pc[8]_i_4_n_0),
        .I0(p_1_in[5])
    );
    LUT1 pc[8]_i_5
    (
        .O(pc[8]_i_5_n_0),
        .I0(p_1_in[4])
    );
    LUT1 pc[8]_i_6
    (
        .O(pc[8]_i_6_n_0),
        .I0(p_1_in[3])
    );
    LUT5 pc[9]_i_2
    (
        .O(pc[9]_i_2_n_0),
        .I0(decodedOpcode_reg_n_0_[0]),
        .I1(decodedOpcode_reg_n_0_[3]),
        .I2(decodedOpcode_reg_n_0_[2]),
        .I3(decodedOpcode_reg_n_0_[4]),
        .I4(decodedOpcode_reg_n_0_[1])
    );
    LUT5 pc[9]_i_3
    (
        .O(pc[9]_i_3_n_0),
        .I0(decodedOpcode_reg_n_0_[0]),
        .I1(decodedOpcode_reg_n_0_[4]),
        .I2(decodedOpcode_reg_n_0_[1]),
        .I3(decodedOpcode_reg_n_0_[2]),
        .I4(decodedOpcode_reg_n_0_[3])
    );
    LUT5 pc[9]_i_4
    (
        .O(pc[9]_i_4_n_0),
        .I0(decodedOpcode_reg_n_0_[0]),
        .I1(decodedOpcode_reg_n_0_[3]),
        .I2(decodedOpcode_reg_n_0_[4]),
        .I3(decodedOpcode_reg_n_0_[1]),
        .I4(decodedOpcode_reg_n_0_[2])
    );
    FDCE pc_reg[0]
    (
        .Q(data0[0]),
        .C(clk_IBUF_BUFG),
        .CE(pc[14]_i_1_n_0),
        .CLR(areset_IBUF),
        .D(pc[0])
    );
    FDCE pc_reg[10]
    (
        .Q(p_1_in[8]),
        .C(clk_IBUF_BUFG),
        .CE(pc[14]_i_1_n_0),
        .CLR(areset_IBUF),
        .D(pc[10])
    );
    FDCE pc_reg[11]
    (
        .Q(p_1_in[9]),
        .C(clk_IBUF_BUFG),
        .CE(pc[14]_i_1_n_0),
        .CLR(areset_IBUF),
        .D(pc[11])
    );
    FDCE pc_reg[12]
    (
        .Q(p_1_in[10]),
        .C(clk_IBUF_BUFG),
        .CE(pc[14]_i_1_n_0),
        .CLR(areset_IBUF),
        .D(pc[12])
    );
    CARRY4 pc_reg[12]_i_2
    (
        .CI(pc_reg[8]_i_2_n_0),
        .CYINIT(<const0>),
        .CO[3:0]({pc_reg[12]_i_2_n_0, pc_reg[12]_i_2_n_1, pc_reg[12]_i_2_n_2, pc_reg[12]_i_2_n_3}),
        .O[3:0]({data2[12], data2[11], data2[10], data2[9]}),
        .DI[3:0]({<const0>, <const0>, <const0>, <const0>}),
        .S[3:0]({pc[12]_i_3_n_0, pc[12]_i_4_n_0, pc[12]_i_5_n_0, pc[12]_i_6_n_0})
    );
    FDCE pc_reg[13]
    (
        .Q(p_1_in[11]),
        .C(clk_IBUF_BUFG),
        .CE(pc[14]_i_1_n_0),
        .CLR(areset_IBUF),
        .D(pc[13])
    );
    FDCE pc_reg[14]
    (
        .Q(p_1_in[12]),
        .C(clk_IBUF_BUFG),
        .CE(pc[14]_i_1_n_0),
        .CLR(areset_IBUF),
        .D(pc[14])
    );
    CARRY4 pc_reg[14]_i_4
    (
        .CI(pc_reg[12]_i_2_n_0),
        .CYINIT(<const0>),
        .CO[3:0]({}),
        .O[3:0]({}),
        .DI[3:0]({<const0>, <const0>, <const0>, <const0>}),
        .S[3:0]({<const0>, <const0>, pc[14]_i_6_n_0, pc[14]_i_7_n_0})
    );
    FDCE pc_reg[1]
    (
        .Q(data0[1]),
        .C(clk_IBUF_BUFG),
        .CE(pc[14]_i_1_n_0),
        .CLR(areset_IBUF),
        .D(pc[1])
    );
    FDCE pc_reg[2]
    (
        .Q(p_1_in[0]),
        .C(clk_IBUF_BUFG),
        .CE(pc[14]_i_1_n_0),
        .CLR(areset_IBUF),
        .D(pc[2])
    );
    FDCE pc_reg[3]
    (
        .Q(p_1_in[1]),
        .C(clk_IBUF_BUFG),
        .CE(pc[14]_i_1_n_0),
        .CLR(areset_IBUF),
        .D(pc[3])
    );
    FDCE pc_reg[4]
    (
        .Q(p_1_in[2]),
        .C(clk_IBUF_BUFG),
        .CE(pc[14]_i_1_n_0),
        .CLR(areset_IBUF),
        .D(pc[4])
    );
    CARRY4 pc_reg[4]_i_2
    (
        .CI(<const0>),
        .CYINIT(data0[0]),
        .CO[3:0]({pc_reg[4]_i_2_n_0, pc_reg[4]_i_2_n_1, pc_reg[4]_i_2_n_2, pc_reg[4]_i_2_n_3}),
        .O[3:0]({data2[4], data2[3], data2[2], data2[1]}),
        .DI[3:0]({<const0>, <const0>, <const0>, <const0>}),
        .S[3:0]({pc[4]_i_3_n_0, pc[4]_i_4_n_0, pc[4]_i_5_n_0, pc[4]_i_6_n_0})
    );
    FDCE pc_reg[5]
    (
        .Q(p_1_in[3]),
        .C(clk_IBUF_BUFG),
        .CE(pc[14]_i_1_n_0),
        .CLR(areset_IBUF),
        .D(pc[5])
    );
    FDCE pc_reg[6]
    (
        .Q(p_1_in[4]),
        .C(clk_IBUF_BUFG),
        .CE(pc[14]_i_1_n_0),
        .CLR(areset_IBUF),
        .D(pc[6])
    );
    FDCE pc_reg[7]
    (
        .Q(p_1_in[5]),
        .C(clk_IBUF_BUFG),
        .CE(pc[14]_i_1_n_0),
        .CLR(areset_IBUF),
        .D(pc[7])
    );
    FDCE pc_reg[8]
    (
        .Q(p_1_in[6]),
        .C(clk_IBUF_BUFG),
        .CE(pc[14]_i_1_n_0),
        .CLR(areset_IBUF),
        .D(pc[8])
    );
    CARRY4 pc_reg[8]_i_2
    (
        .CI(pc_reg[4]_i_2_n_0),
        .CYINIT(<const0>),
        .CO[3:0]({pc_reg[8]_i_2_n_0, pc_reg[8]_i_2_n_1, pc_reg[8]_i_2_n_2, pc_reg[8]_i_2_n_3}),
        .O[3:0]({data2[8], data2[7], data2[6], data2[5]}),
        .DI[3:0]({<const0>, <const0>, <const0>, <const0>}),
        .S[3:0]({pc[8]_i_3_n_0, pc[8]_i_4_n_0, pc[8]_i_5_n_0, pc[8]_i_6_n_0})
    );
    FDCE pc_reg[9]
    (
        .Q(p_1_in[7]),
        .C(clk_IBUF_BUFG),
        .CE(pc[14]_i_1_n_0),
        .CLR(areset_IBUF),
        .D(pc[9])
    );
    LUT1 sp[10]_i_10
    (
        .O(sp[10]_i_10_n_0),
        .I0(sp_reg_n_0_[9])
    );
    LUT1 sp[10]_i_11
    (
        .O(sp[10]_i_11_n_0),
        .I0(sp_reg_n_0_[8])
    );
    LUT1 sp[10]_i_12
    (
        .O(sp[10]_i_12_n_0),
        .I0(sp_reg_n_0_[7])
    );
    LUT1 sp[10]_i_5
    (
        .O(sp[10]_i_5_n_0),
        .I0(sp_reg_n_0_[10])
    );
    LUT1 sp[10]_i_6
    (
        .O(sp[10]_i_6_n_0),
        .I0(sp_reg_n_0_[9])
    );
    LUT1 sp[10]_i_7
    (
        .O(sp[10]_i_7_n_0),
        .I0(sp_reg_n_0_[8])
    );
    LUT1 sp[10]_i_8
    (
        .O(sp[10]_i_8_n_0),
        .I0(sp_reg_n_0_[7])
    );
    LUT1 sp[10]_i_9
    (
        .O(sp[10]_i_9_n_0),
        .I0(sp_reg_n_0_[10])
    );
    LUT5 sp[14]_i_1
    (
        .O(sp[14]_i_1_n_0),
        .I0(g0_b0__0_n_0),
        .I1(FSM_sequential_state_reg_n_0_[0]),
        .I2(FSM_sequential_state_reg_n_0_[2]),
        .I3(FSM_sequential_state_reg_n_0_[1]),
        .I4(FSM_sequential_state_reg_n_0_[3])
    );
    LUT1 sp[14]_i_10
    (
        .O(sp[14]_i_10_n_0),
        .I0(sp_reg_n_0_[13])
    );
    LUT1 sp[14]_i_11
    (
        .O(sp[14]_i_11_n_0),
        .I0(sp_reg_n_0_[12])
    );
    LUT1 sp[14]_i_12
    (
        .O(sp[14]_i_12_n_0),
        .I0(sp_reg_n_0_[11])
    );
    LUT1 sp[14]_i_13
    (
        .O(sp[14]_i_13_n_0),
        .I0(sp_reg_n_0_[14])
    );
    LUT1 sp[14]_i_14
    (
        .O(sp[14]_i_14_n_0),
        .I0(sp_reg_n_0_[13])
    );
    LUT1 sp[14]_i_15
    (
        .O(sp[14]_i_15_n_0),
        .I0(sp_reg_n_0_[12])
    );
    LUT1 sp[14]_i_16
    (
        .O(sp[14]_i_16_n_0),
        .I0(sp_reg_n_0_[11])
    );
    LUT4 sp[14]_i_4
    (
        .O(sp[14]_i_4_n_0),
        .I0(decodedOpcode_reg_n_0_[2]),
        .I1(decodedOpcode_reg_n_0_[0]),
        .I2(decodedOpcode_reg_n_0_[1]),
        .I3(decodedOpcode_reg_n_0_[3])
    );
    LUT6 sp[14]_i_6
    (
        .O(sp[14]_i_6_n_0),
        .I0(decodedOpcode_reg_n_0_[2]),
        .I1(decodedOpcode_reg_n_0_[3]),
        .I2(decodedOpcode_reg_n_0_[1]),
        .I3(decodedOpcode_reg_n_0_[0]),
        .I4(idim_flag),
        .I5(decodedOpcode_reg_n_0_[4])
    );
    LUT4 sp[14]_i_8
    (
        .O(sp[14]_i_8_n_0),
        .I0(decodedOpcode_reg_n_0_[0]),
        .I1(decodedOpcode_reg_n_0_[1]),
        .I2(decodedOpcode_reg_n_0_[3]),
        .I3(decodedOpcode_reg_n_0_[4])
    );
    LUT1 sp[14]_i_9
    (
        .O(sp[14]_i_9_n_0),
        .I0(sp_reg_n_0_[14])
    );
    LUT5 sp[2]_i_2
    (
        .O(sp[2]_i_2_n_0),
        .I0(decodedOpcode_reg_n_0_[4]),
        .I1(decodedOpcode_reg_n_0_[3]),
        .I2(decodedOpcode_reg_n_0_[1]),
        .I3(decodedOpcode_reg_n_0_[0]),
        .I4(idim_flag)
    );
    LUT1 sp[6]_i_10
    (
        .O(sp[6]_i_10_n_0),
        .I0(sp_reg_n_0_[5])
    );
    LUT1 sp[6]_i_11
    (
        .O(sp[6]_i_11_n_0),
        .I0(sp_reg_n_0_[4])
    );
    LUT1 sp[6]_i_12
    (
        .O(sp[6]_i_12_n_0),
        .I0(sp_reg_n_0_[3])
    );
    LUT1 sp[6]_i_5
    (
        .O(sp[6]_i_5_n_0),
        .I0(sp_reg_n_0_[6])
    );
    LUT1 sp[6]_i_6
    (
        .O(sp[6]_i_6_n_0),
        .I0(sp_reg_n_0_[5])
    );
    LUT1 sp[6]_i_7
    (
        .O(sp[6]_i_7_n_0),
        .I0(sp_reg_n_0_[4])
    );
    LUT1 sp[6]_i_8
    (
        .O(sp[6]_i_8_n_0),
        .I0(sp_reg_n_0_[3])
    );
    LUT1 sp[6]_i_9
    (
        .O(sp[6]_i_9_n_0),
        .I0(sp_reg_n_0_[6])
    );
    FDPE sp_reg[10]
    (
        .Q(sp_reg_n_0_[10]),
        .C(clk_IBUF_BUFG),
        .CE(sp[14]_i_1_n_0),
        .D(sp[10]),
        .PRE(areset_IBUF)
    );
    CARRY4 sp_reg[10]_i_3
    (
        .CI(sp_reg[6]_i_3_n_0),
        .CYINIT(<const0>),
        .CO[3:0]({sp_reg[10]_i_3_n_0, sp_reg[10]_i_3_n_1, sp_reg[10]_i_3_n_2, sp_reg[10]_i_3_n_3}),
        .O[3:0]({sp_reg[10]_i_3_n_4, sp_reg[10]_i_3_n_5, sp_reg[10]_i_3_n_6, sp_reg[10]_i_3_n_7}),
        .DI[3:0]({<const0>, <const0>, <const0>, <const0>}),
        .S[3:0]({sp[10]_i_5_n_0, sp[10]_i_6_n_0, sp[10]_i_7_n_0, sp[10]_i_8_n_0})
    );
    CARRY4 sp_reg[10]_i_4
    (
        .CI(sp_reg[6]_i_4_n_0),
        .CYINIT(<const0>),
        .CO[3:0]({sp_reg[10]_i_4_n_0, sp_reg[10]_i_4_n_1, sp_reg[10]_i_4_n_2, sp_reg[10]_i_4_n_3}),
        .O[3:0]({sp_reg[10]_i_4_n_4, sp_reg[10]_i_4_n_5, sp_reg[10]_i_4_n_6, sp_reg[10]_i_4_n_7}),
        .DI[3:0]({sp_reg_n_0_[10], sp_reg_n_0_[9], sp_reg_n_0_[8], sp_reg_n_0_[7]}),
        .S[3:0]({sp[10]_i_9_n_0, sp[10]_i_10_n_0, sp[10]_i_11_n_0, sp[10]_i_12_n_0})
    );
    FDPE sp_reg[11]
    (
        .Q(sp_reg_n_0_[11]),
        .C(clk_IBUF_BUFG),
        .CE(sp[14]_i_1_n_0),
        .D(sp[11]),
        .PRE(areset_IBUF)
    );
    FDPE sp_reg[12]
    (
        .Q(sp_reg_n_0_[12]),
        .C(clk_IBUF_BUFG),
        .CE(sp[14]_i_1_n_0),
        .D(sp[12]),
        .PRE(areset_IBUF)
    );
    FDPE sp_reg[13]
    (
        .Q(sp_reg_n_0_[13]),
        .C(clk_IBUF_BUFG),
        .CE(sp[14]_i_1_n_0),
        .D(sp[13]),
        .PRE(areset_IBUF)
    );
    FDPE sp_reg[14]
    (
        .Q(sp_reg_n_0_[14]),
        .C(clk_IBUF_BUFG),
        .CE(sp[14]_i_1_n_0),
        .D(sp[14]),
        .PRE(areset_IBUF)
    );
    CARRY4 sp_reg[14]_i_5
    (
        .CI(sp_reg[10]_i_3_n_0),
        .CYINIT(<const0>),
        .CO[3:0]({}),
        .O[3:0]({sp_reg[14]_i_5_n_4, sp_reg[14]_i_5_n_5, sp_reg[14]_i_5_n_6, sp_reg[14]_i_5_n_7}),
        .DI[3:0]({<const0>, <const0>, <const0>, <const0>}),
        .S[3:0]({sp[14]_i_9_n_0, sp[14]_i_10_n_0, sp[14]_i_11_n_0, sp[14]_i_12_n_0})
    );
    CARRY4 sp_reg[14]_i_7
    (
        .CI(sp_reg[10]_i_4_n_0),
        .CYINIT(<const0>),
        .CO[3:0]({}),
        .O[3:0]({sp_reg[14]_i_7_n_4, sp_reg[14]_i_7_n_5, sp_reg[14]_i_7_n_6, sp_reg[14]_i_7_n_7}),
        .DI[3:0]({<const0>, sp_reg_n_0_[13], sp_reg_n_0_[12], sp_reg_n_0_[11]}),
        .S[3:0]({sp[14]_i_13_n_0, sp[14]_i_14_n_0, sp[14]_i_15_n_0, sp[14]_i_16_n_0})
    );
    FDCE sp_reg[2]
    (
        .Q(sp_reg_n_0_[2]),
        .C(clk_IBUF_BUFG),
        .CE(sp[14]_i_1_n_0),
        .CLR(areset_IBUF),
        .D(sp[2])
    );
    FDPE sp_reg[3]
    (
        .Q(sp_reg_n_0_[3]),
        .C(clk_IBUF_BUFG),
        .CE(sp[14]_i_1_n_0),
        .D(sp[3]),
        .PRE(areset_IBUF)
    );
    FDPE sp_reg[4]
    (
        .Q(sp_reg_n_0_[4]),
        .C(clk_IBUF_BUFG),
        .CE(sp[14]_i_1_n_0),
        .D(sp[4]),
        .PRE(areset_IBUF)
    );
    FDPE sp_reg[5]
    (
        .Q(sp_reg_n_0_[5]),
        .C(clk_IBUF_BUFG),
        .CE(sp[14]_i_1_n_0),
        .D(sp[5]),
        .PRE(areset_IBUF)
    );
    FDPE sp_reg[6]
    (
        .Q(sp_reg_n_0_[6]),
        .C(clk_IBUF_BUFG),
        .CE(sp[14]_i_1_n_0),
        .D(sp[6]),
        .PRE(areset_IBUF)
    );
    CARRY4 sp_reg[6]_i_3
    (
        .CI(<const0>),
        .CYINIT(sp_reg_n_0_[2]),
        .CO[3:0]({sp_reg[6]_i_3_n_0, sp_reg[6]_i_3_n_1, sp_reg[6]_i_3_n_2, sp_reg[6]_i_3_n_3}),
        .O[3:0]({sp_reg[6]_i_3_n_4, sp_reg[6]_i_3_n_5, sp_reg[6]_i_3_n_6, sp_reg[6]_i_3_n_7}),
        .DI[3:0]({<const0>, <const0>, <const0>, <const0>}),
        .S[3:0]({sp[6]_i_5_n_0, sp[6]_i_6_n_0, sp[6]_i_7_n_0, sp[6]_i_8_n_0})
    );
    CARRY4 sp_reg[6]_i_4
    (
        .CI(<const0>),
        .CYINIT(sp_reg_n_0_[2]),
        .CO[3:0]({sp_reg[6]_i_4_n_0, sp_reg[6]_i_4_n_1, sp_reg[6]_i_4_n_2, sp_reg[6]_i_4_n_3}),
        .O[3:0]({sp_reg[6]_i_4_n_4, sp_reg[6]_i_4_n_5, sp_reg[6]_i_4_n_6, sp_reg[6]_i_4_n_7}),
        .DI[3:0]({sp_reg_n_0_[6], sp_reg_n_0_[5], sp_reg_n_0_[4], sp_reg_n_0_[3]}),
        .S[3:0]({sp[6]_i_9_n_0, sp[6]_i_10_n_0, sp[6]_i_11_n_0, sp[6]_i_12_n_0})
    );
    FDPE sp_reg[7]
    (
        .Q(sp_reg_n_0_[7]),
        .C(clk_IBUF_BUFG),
        .CE(sp[14]_i_1_n_0),
        .D(sp[7]),
        .PRE(areset_IBUF)
    );
    FDPE sp_reg[8]
    (
        .Q(sp_reg_n_0_[8]),
        .C(clk_IBUF_BUFG),
        .CE(sp[14]_i_1_n_0),
        .D(sp[8]),
        .PRE(areset_IBUF)
    );
    FDPE sp_reg[9]
    (
        .Q(sp_reg_n_0_[9]),
        .C(clk_IBUF_BUFG),
        .CE(sp[14]_i_1_n_0),
        .D(sp[9]),
        .PRE(areset_IBUF)
    );
endmodule

module LUT6
(
    O,
    I0,
    I1,
    I2,
    I3,
    I4,
    I5
);

    output O;
    input I0;
    input I1;
    input I2;
    input I3;
    input I4;
    input I5;


endmodule

module LUT2
(
    O,
    I0,
    I1
);

    output O;
    input I0;
    input I1;


endmodule

module LUT4
(
    O,
    I0,
    I1,
    I2,
    I3
);

    output O;
    input I0;
    input I1;
    input I2;
    input I3;


endmodule

module LUT5
(
    O,
    I0,
    I1,
    I2,
    I3,
    I4
);

    output O;
    input I0;
    input I1;
    input I2;
    input I3;
    input I4;


endmodule

module FDCE
(
    Q,
    C,
    CE,
    CLR,
    D
);

    output Q;
    input C;
    input CE;
    input CLR;
    input D;


endmodule

module GND
(
    G
);

    output G;


endmodule

module VCC
(
    P
);

    output P;


endmodule

module IBUF
(
    O,
    I
);

    output O;
    input I;


endmodule

module OBUF
(
    O,
    I
);

    output O;
    input I;


endmodule

module BUFG
(
    O,
    I
);

    output O;
    input I;


endmodule

module LUT3
(
    O,
    I0,
    I1,
    I2
);

    output O;
    input I0;
    input I1;
    input I2;


endmodule

module FDRE
(
    Q,
    C,
    CE,
    D,
    R
);

    output Q;
    input C;
    input CE;
    input D;
    input R;


endmodule

module LUT1
(
    O,
    I0
);

    output O;
    input I0;


endmodule

module CARRY4
(
    CI,
    CYINIT,
    CO[3:0],
    O[3:0],
    DI[3:0],
    S[3:0]
);

    input CI;
    input CYINIT;
    output [3:0]CO[3:0];
    output [3:0]O[3:0];
    input [3:0]DI[3:0];
    input [3:0]S[3:0];


endmodule

module dualport_ram
(
    .FSM_sequential_state_reg[0]({FSM_sequential_state_reg[0]}),
    .FSM_sequential_state_reg[1]({FSM_sequential_state_reg[1]}),
    FSM_sequential_state_reg[1]_0,
    .FSM_sequential_state_reg[2]({FSM_sequential_state_reg[2]}),
    .FSM_sequential_state_reg[3]({FSM_sequential_state_reg[3]}),
    clk_IBUF_BUFG,
    .decodedOpcode_reg[0]({decodedOpcode_reg[0]}),
    decodedOpcode_reg[0]_0,
    decodedOpcode_reg[0]_1,
    decodedOpcode_reg[0]_2,
    decodedOpcode_reg[0]_3,
    decodedOpcode_reg[0]_4,
    .decodedOpcode_reg[1]({decodedOpcode_reg[1]}),
    .decodedOpcode_reg[2]({decodedOpcode_reg[2]}),
    decodedOpcode_reg[2]_0,
    decodedOpcode_reg[2]_1,
    decodedOpcode_reg[2]_10,
    decodedOpcode_reg[2]_11,
    decodedOpcode_reg[2]_12,
    decodedOpcode_reg[2]_13,
    decodedOpcode_reg[2]_14,
    decodedOpcode_reg[2]_15,
    decodedOpcode_reg[2]_16,
    decodedOpcode_reg[2]_17,
    decodedOpcode_reg[2]_2,
    decodedOpcode_reg[2]_3,
    decodedOpcode_reg[2]_4,
    decodedOpcode_reg[2]_5,
    decodedOpcode_reg[2]_6,
    decodedOpcode_reg[2]_7,
    decodedOpcode_reg[2]_8,
    decodedOpcode_reg[2]_9,
    .decodedOpcode_reg[3]({decodedOpcode_reg[3]}),
    decodedOpcode_reg[3]_0,
    decodedOpcode_reg[3]_1,
    decodedOpcode_reg[3]_10,
    decodedOpcode_reg[3]_11,
    decodedOpcode_reg[3]_12,
    decodedOpcode_reg[3]_2,
    decodedOpcode_reg[3]_3,
    decodedOpcode_reg[3]_4,
    decodedOpcode_reg[3]_5,
    decodedOpcode_reg[3]_6,
    decodedOpcode_reg[3]_7,
    decodedOpcode_reg[3]_8,
    decodedOpcode_reg[3]_9,
    decodedOpcode_reg[4]_0,
    decodedOpcode_reg[4]_1,
    idim_flag,
    inInterrupt_reg,
    in_mem_busy_IBUF,
    memAWriteEnable,
    memBWriteEnable,
    .opcode_reg[0]({opcode_reg[0]}),
    opcode_reg[0]_0,
    opcode_reg[0]_1,
    .opcode_reg[1]({opcode_reg[1]}),
    opcode_reg[1]_0,
    .opcode_reg[2]({opcode_reg[2]}),
    .opcode_reg[3]({opcode_reg[3]}),
    .opcode_reg[4]({opcode_reg[4]}),
    .opcode_reg[5]({opcode_reg[5]}),
    .opcode_reg[6]({opcode_reg[6]}),
    out_mem_readEnable_reg,
    .pc_reg[10]({pc_reg[10]}),
    .pc_reg[11]({pc_reg[11]}),
    .pc_reg[12]({pc_reg[12]}),
    .pc_reg[13]({pc_reg[13]}),
    pc_reg[14]_0,
    .pc_reg[2]({pc_reg[2]}),
    .pc_reg[3]({pc_reg[3]}),
    .pc_reg[4]({pc_reg[4]}),
    .pc_reg[5]({pc_reg[5]}),
    .pc_reg[6]({pc_reg[6]}),
    .pc_reg[7]({pc_reg[7]}),
    .pc_reg[8]({pc_reg[8]}),
    .pc_reg[9]({pc_reg[9]}),
    .D[2:0]({D[2], D[1], D[0]}),
    .O[3:0]({O[3], O[2], O[1], O[0]}),
    .Q[4:0]({Q[4], Q[3], Q[2], Q[1], Q[0]}),
    .data2[11:0]({data2[11], data2[10], data2[9], data2[8], data2[7], data2[6], data2[5], data2[4], data2[3], data2[2], data2[1], data2[0]}),
    .decodedOpcode_reg[4][4:0]({decodedOpcode_reg[4][4], decodedOpcode_reg[4][3], decodedOpcode_reg[4][2], decodedOpcode_reg[4][1], decodedOpcode_reg[4][0]}),
    .memAAddr_reg[14][12:0]({memAAddr_reg[14][12], memAAddr_reg[14][11], memAAddr_reg[14][10], memAAddr_reg[14][9], memAAddr_reg[14][8], memAAddr_reg[14][7], memAAddr_reg[14][6], memAAddr_reg[14][5], memAAddr_reg[14][4], memAAddr_reg[14][3], memAAddr_reg[14][2], memAAddr_reg[14][1], memAAddr_reg[14][0]}),
    .memAAddr_reg[14]_0[12:0]({memAAddr_reg[14]_0[12], memAAddr_reg[14]_0[11], memAAddr_reg[14]_0[10], memAAddr_reg[14]_0[9], memAAddr_reg[14]_0[8], memAAddr_reg[14]_0[7], memAAddr_reg[14]_0[6], memAAddr_reg[14]_0[5], memAAddr_reg[14]_0[4], memAAddr_reg[14]_0[3], memAAddr_reg[14]_0[2], memAAddr_reg[14]_0[1], memAAddr_reg[14]_0[0]}),
    .memARead[31:0]({memARead[31], memARead[30], memARead[29], memARead[28], memARead[27], memARead[26], memARead[25], memARead[24], memARead[23], memARead[22], memARead[21], memARead[20], memARead[19], memARead[18], memARead[17], memARead[16], memARead[15], memARead[14], memARead[13], memARead[12], memARead[11], memARead[10], memARead[9], memARead[8], memARead[7], memARead[6], memARead[5], memARead[4], memARead[3], memARead[2], memARead[1], memARead[0]}),
    .memAWrite_reg[31][31:0]({memAWrite_reg[31][31], memAWrite_reg[31][30], memAWrite_reg[31][29], memAWrite_reg[31][28], memAWrite_reg[31][27], memAWrite_reg[31][26], memAWrite_reg[31][25], memAWrite_reg[31][24], memAWrite_reg[31][23], memAWrite_reg[31][22], memAWrite_reg[31][21], memAWrite_reg[31][20], memAWrite_reg[31][19], memAWrite_reg[31][18], memAWrite_reg[31][17], memAWrite_reg[31][16], memAWrite_reg[31][15], memAWrite_reg[31][14], memAWrite_reg[31][13], memAWrite_reg[31][12], memAWrite_reg[31][11], memAWrite_reg[31][10], memAWrite_reg[31][9], memAWrite_reg[31][8], memAWrite_reg[31][7], memAWrite_reg[31][6], memAWrite_reg[31][5], memAWrite_reg[31][4], memAWrite_reg[31][3], memAWrite_reg[31][2], memAWrite_reg[31][1], memAWrite_reg[31][0]}),
    .memAWrite_reg[31]_0[31:0]({memAWrite_reg[31]_0[31], memAWrite_reg[31]_0[30], memAWrite_reg[31]_0[29], memAWrite_reg[31]_0[28], memAWrite_reg[31]_0[27], memAWrite_reg[31]_0[26], memAWrite_reg[31]_0[25], memAWrite_reg[31]_0[24], memAWrite_reg[31]_0[23], memAWrite_reg[31]_0[22], memAWrite_reg[31]_0[21], memAWrite_reg[31]_0[20], memAWrite_reg[31]_0[19], memAWrite_reg[31]_0[18], memAWrite_reg[31]_0[17], memAWrite_reg[31]_0[16], memAWrite_reg[31]_0[15], memAWrite_reg[31]_0[14], memAWrite_reg[31]_0[13], memAWrite_reg[31]_0[12], memAWrite_reg[31]_0[11], memAWrite_reg[31]_0[10], memAWrite_reg[31]_0[9], memAWrite_reg[31]_0[8], memAWrite_reg[31]_0[7], memAWrite_reg[31]_0[6], memAWrite_reg[31]_0[5], memAWrite_reg[31]_0[4], memAWrite_reg[31]_0[3], memAWrite_reg[31]_0[2], memAWrite_reg[31]_0[1], memAWrite_reg[31]_0[0]}),
    .memBAddr_reg[14][12:0]({memBAddr_reg[14][12], memBAddr_reg[14][11], memBAddr_reg[14][10], memBAddr_reg[14][9], memBAddr_reg[14][8], memBAddr_reg[14][7], memBAddr_reg[14][6], memBAddr_reg[14][5], memBAddr_reg[14][4], memBAddr_reg[14][3], memBAddr_reg[14][2], memBAddr_reg[14][1], memBAddr_reg[14][0]}),
    .memBRead[31:0]({memBRead[31], memBRead[30], memBRead[29], memBRead[28], memBRead[27], memBRead[26], memBRead[25], memBRead[24], memBRead[23], memBRead[22], memBRead[21], memBRead[20], memBRead[19], memBRead[18], memBRead[17], memBRead[16], memBRead[15], memBRead[14], memBRead[13], memBRead[12], memBRead[11], memBRead[10], memBRead[9], memBRead[8], memBRead[7], memBRead[6], memBRead[5], memBRead[4], memBRead[3], memBRead[2], memBRead[1], memBRead[0]}),
    .memBWrite_reg[31][31:0]({memBWrite_reg[31][31], memBWrite_reg[31][30], memBWrite_reg[31][29], memBWrite_reg[31][28], memBWrite_reg[31][27], memBWrite_reg[31][26], memBWrite_reg[31][25], memBWrite_reg[31][24], memBWrite_reg[31][23], memBWrite_reg[31][22], memBWrite_reg[31][21], memBWrite_reg[31][20], memBWrite_reg[31][19], memBWrite_reg[31][18], memBWrite_reg[31][17], memBWrite_reg[31][16], memBWrite_reg[31][15], memBWrite_reg[31][14], memBWrite_reg[31][13], memBWrite_reg[31][12], memBWrite_reg[31][11], memBWrite_reg[31][10], memBWrite_reg[31][9], memBWrite_reg[31][8], memBWrite_reg[31][7], memBWrite_reg[31][6], memBWrite_reg[31][5], memBWrite_reg[31][4], memBWrite_reg[31][3], memBWrite_reg[31][2], memBWrite_reg[31][1], memBWrite_reg[31][0]}),
    .mem_read_IBUF[31:0]({mem_read_IBUF[31], mem_read_IBUF[30], mem_read_IBUF[29], mem_read_IBUF[28], mem_read_IBUF[27], mem_read_IBUF[26], mem_read_IBUF[25], mem_read_IBUF[24], mem_read_IBUF[23], mem_read_IBUF[22], mem_read_IBUF[21], mem_read_IBUF[20], mem_read_IBUF[19], mem_read_IBUF[18], mem_read_IBUF[17], mem_read_IBUF[16], mem_read_IBUF[15], mem_read_IBUF[14], mem_read_IBUF[13], mem_read_IBUF[12], mem_read_IBUF[11], mem_read_IBUF[10], mem_read_IBUF[9], mem_read_IBUF[8], mem_read_IBUF[7], mem_read_IBUF[6], mem_read_IBUF[5], mem_read_IBUF[4], mem_read_IBUF[3], mem_read_IBUF[2], mem_read_IBUF[1], mem_read_IBUF[0]}),
    .opcode_reg[6]_0[4:0]({opcode_reg[6]_0[4], opcode_reg[6]_0[3], opcode_reg[6]_0[2], opcode_reg[6]_0[1], opcode_reg[6]_0[0]}),
    .out[3:0]({out[3], out[2], out[1], out[0]}),
    .pc_reg[14][14:0]({pc_reg[14][14], pc_reg[14][13], pc_reg[14][12], pc_reg[14][11], pc_reg[14][10], pc_reg[14][9], pc_reg[14][8], pc_reg[14][7], pc_reg[14][6], pc_reg[14][5], pc_reg[14][4], pc_reg[14][3], pc_reg[14][2], pc_reg[14][1], pc_reg[14][0]}),
    .pc_reg[14]_1[13:0]({pc_reg[14]_1[13], pc_reg[14]_1[12], pc_reg[14]_1[11], pc_reg[14]_1[10], pc_reg[14]_1[9], pc_reg[14]_1[8], pc_reg[14]_1[7], pc_reg[14]_1[6], pc_reg[14]_1[5], pc_reg[14]_1[4], pc_reg[14]_1[3], pc_reg[14]_1[2], pc_reg[14]_1[1], pc_reg[14]_1[0]}),
    .pc_reg[1][1:0]({pc_reg[1][1], pc_reg[1][0]}),
    .sp_reg[10][3:0]({sp_reg[10][3], sp_reg[10][2], sp_reg[10][1], sp_reg[10][0]}),
    .sp_reg[14][12:0]({sp_reg[14][12], sp_reg[14][11], sp_reg[14][10], sp_reg[14][9], sp_reg[14][8], sp_reg[14][7], sp_reg[14][6], sp_reg[14][5], sp_reg[14][4], sp_reg[14][3], sp_reg[14][2], sp_reg[14][1], sp_reg[14][0]}),
    .sp_reg[14]_0[12:0]({sp_reg[14]_0[12], sp_reg[14]_0[11], sp_reg[14]_0[10], sp_reg[14]_0[9], sp_reg[14]_0[8], sp_reg[14]_0[7], sp_reg[14]_0[6], sp_reg[14]_0[5], sp_reg[14]_0[4], sp_reg[14]_0[3], sp_reg[14]_0[2], sp_reg[14]_0[1], sp_reg[14]_0[0]}),
    .sp_reg[2][3:0]({sp_reg[2][3], sp_reg[2][2], sp_reg[2][1], sp_reg[2][0]})
);

    input [3:0]FSM_sequential_state_reg;
    input [3:0]FSM_sequential_state_reg;
    input FSM_sequential_state_reg[1]_0;
    input [3:0]FSM_sequential_state_reg;
    input [3:0]FSM_sequential_state_reg;
    input clk_IBUF_BUFG;
    input [3:0]decodedOpcode_reg;
    input decodedOpcode_reg[0]_0;
    input decodedOpcode_reg[0]_1;
    input decodedOpcode_reg[0]_2;
    input decodedOpcode_reg[0]_3;
    input decodedOpcode_reg[0]_4;
    input [3:0]decodedOpcode_reg;
    input [3:0]decodedOpcode_reg;
    input decodedOpcode_reg[2]_0;
    input decodedOpcode_reg[2]_1;
    input decodedOpcode_reg[2]_10;
    input decodedOpcode_reg[2]_11;
    input decodedOpcode_reg[2]_12;
    input decodedOpcode_reg[2]_13;
    input decodedOpcode_reg[2]_14;
    input decodedOpcode_reg[2]_15;
    input decodedOpcode_reg[2]_16;
    input decodedOpcode_reg[2]_17;
    input decodedOpcode_reg[2]_2;
    input decodedOpcode_reg[2]_3;
    input decodedOpcode_reg[2]_4;
    input decodedOpcode_reg[2]_5;
    input decodedOpcode_reg[2]_6;
    input decodedOpcode_reg[2]_7;
    input decodedOpcode_reg[2]_8;
    input decodedOpcode_reg[2]_9;
    input [3:0]decodedOpcode_reg;
    input decodedOpcode_reg[3]_0;
    input decodedOpcode_reg[3]_1;
    input decodedOpcode_reg[3]_10;
    input decodedOpcode_reg[3]_11;
    input decodedOpcode_reg[3]_12;
    input decodedOpcode_reg[3]_2;
    input decodedOpcode_reg[3]_3;
    input decodedOpcode_reg[3]_4;
    input decodedOpcode_reg[3]_5;
    input decodedOpcode_reg[3]_6;
    input decodedOpcode_reg[3]_7;
    input decodedOpcode_reg[3]_8;
    input decodedOpcode_reg[3]_9;
    input decodedOpcode_reg[4]_0;
    input decodedOpcode_reg[4]_1;
    input idim_flag;
    input inInterrupt_reg;
    input in_mem_busy_IBUF;
    input memAWriteEnable;
    input memBWriteEnable;
    output [6:0]opcode_reg;
    input opcode_reg[0]_0;
    input opcode_reg[0]_1;
    output [6:0]opcode_reg;
    input opcode_reg[1]_0;
    output [6:0]opcode_reg;
    output [6:0]opcode_reg;
    output [6:0]opcode_reg;
    output [6:0]opcode_reg;
    output [6:0]opcode_reg;
    output out_mem_readEnable_reg;
    input [13:2]pc_reg;
    input [13:2]pc_reg;
    input [13:2]pc_reg;
    input [13:2]pc_reg;
    input pc_reg[14]_0;
    input [13:2]pc_reg;
    input [13:2]pc_reg;
    input [13:2]pc_reg;
    input [13:2]pc_reg;
    input [13:2]pc_reg;
    input [13:2]pc_reg;
    input [13:2]pc_reg;
    input [13:2]pc_reg;
    output [2:0]D;
    input [3:0]O;
    input [4:0]Q;
    input [11:0]data2;
    output [4:0]decodedOpcode_reg[4];
    output [12:0]memAAddr_reg[14];
    input [12:0]memAAddr_reg[14]_0;
    output [31:0]memARead;
    output [31:0]memAWrite_reg[31];
    input [31:0]memAWrite_reg[31]_0;
    input [12:0]memBAddr_reg[14];
    output [31:0]memBRead;
    input [31:0]memBWrite_reg[31];
    input [31:0]mem_read_IBUF;
    input [4:0]opcode_reg[6]_0;
    input [3:0]out;
    output [14:0]pc_reg[14];
    input [13:0]pc_reg[14]_1;
    input [1:0]pc_reg[1];
    input [3:0]sp_reg[10];
    output [12:0]sp_reg[14];
    input [12:0]sp_reg[14]_0;
    input [3:0]sp_reg[2];

    wire <const0>;
    wire <const1>;
    wire [2:0]D;
    wire FSM_sequential_state[1]_i_2_n_0;
    wire FSM_sequential_state[2]_i_2_n_0;
    wire FSM_sequential_state[3]_i_4_n_0;
    wire [3:0]FSM_sequential_state_reg;
    wire FSM_sequential_state_reg[1]_0;
    wire [3:0]O;
    wire [4:0]Q;
    wire clk_IBUF_BUFG;
    wire [11:0]data2;
    wire decodedOpcode[0]_i_2_n_0;
    wire decodedOpcode[1]_i_2_n_0;
    wire decodedOpcode[2]_i_2_n_0;
    wire decodedOpcode[2]_i_3_n_0;
    wire decodedOpcode[2]_i_4_n_0;
    wire decodedOpcode[3]_i_2_n_0;
    wire decodedOpcode[3]_i_3_n_0;
    wire decodedOpcode[4]_i_3_n_0;
    wire decodedOpcode[4]_i_4_n_0;
    wire [3:0]decodedOpcode_reg;
    wire decodedOpcode_reg[0]_0;
    wire decodedOpcode_reg[0]_1;
    wire decodedOpcode_reg[0]_2;
    wire decodedOpcode_reg[0]_3;
    wire decodedOpcode_reg[0]_4;
    wire decodedOpcode_reg[2]_0;
    wire decodedOpcode_reg[2]_1;
    wire decodedOpcode_reg[2]_10;
    wire decodedOpcode_reg[2]_11;
    wire decodedOpcode_reg[2]_12;
    wire decodedOpcode_reg[2]_13;
    wire decodedOpcode_reg[2]_14;
    wire decodedOpcode_reg[2]_15;
    wire decodedOpcode_reg[2]_16;
    wire decodedOpcode_reg[2]_17;
    wire decodedOpcode_reg[2]_2;
    wire decodedOpcode_reg[2]_3;
    wire decodedOpcode_reg[2]_4;
    wire decodedOpcode_reg[2]_5;
    wire decodedOpcode_reg[2]_6;
    wire decodedOpcode_reg[2]_7;
    wire decodedOpcode_reg[2]_8;
    wire decodedOpcode_reg[2]_9;
    wire decodedOpcode_reg[3]_0;
    wire decodedOpcode_reg[3]_1;
    wire decodedOpcode_reg[3]_10;
    wire decodedOpcode_reg[3]_11;
    wire decodedOpcode_reg[3]_12;
    wire decodedOpcode_reg[3]_2;
    wire decodedOpcode_reg[3]_3;
    wire decodedOpcode_reg[3]_4;
    wire decodedOpcode_reg[3]_5;
    wire decodedOpcode_reg[3]_6;
    wire decodedOpcode_reg[3]_7;
    wire decodedOpcode_reg[3]_8;
    wire decodedOpcode_reg[3]_9;
    wire [4:0]decodedOpcode_reg[4];
    wire decodedOpcode_reg[4]_0;
    wire decodedOpcode_reg[4]_1;
    wire idim_flag;
    wire inInterrupt_reg;
    wire in_mem_busy_IBUF;
    wire memAAddr[10]_i_2_n_0;
    wire memAAddr[10]_i_3_n_0;
    wire memAAddr[11]_i_2_n_0;
    wire memAAddr[11]_i_3_n_0;
    wire memAAddr[12]_i_2_n_0;
    wire memAAddr[12]_i_3_n_0;
    wire memAAddr[13]_i_2_n_0;
    wire memAAddr[13]_i_3_n_0;
    wire memAAddr[14]_i_2_n_0;
    wire memAAddr[14]_i_3_n_0;
    wire memAAddr[2]_i_2_n_0;
    wire memAAddr[3]_i_2_n_0;
    wire memAAddr[3]_i_3_n_0;
    wire memAAddr[4]_i_2_n_0;
    wire memAAddr[4]_i_3_n_0;
    wire memAAddr[5]_i_2_n_0;
    wire memAAddr[5]_i_3_n_0;
    wire memAAddr[6]_i_2_n_0;
    wire memAAddr[6]_i_3_n_0;
    wire memAAddr[7]_i_2_n_0;
    wire memAAddr[7]_i_3_n_0;
    wire memAAddr[8]_i_2_n_0;
    wire memAAddr[8]_i_3_n_0;
    wire memAAddr[9]_i_2_n_0;
    wire memAAddr[9]_i_3_n_0;
    wire [12:0]memAAddr_reg[14];
    wire [12:0]memAAddr_reg[14]_0;
    wire [31:0]memARead;
    wire memAWriteEnable;
    wire memAWrite[0]_i_2_n_0;
    wire memAWrite[0]_i_3_n_0;
    wire memAWrite[0]_i_5_n_0;
    wire memAWrite[10]_i_2_n_0;
    wire memAWrite[10]_i_3_n_0;
    wire memAWrite[10]_i_5_n_0;
    wire memAWrite[10]_i_6_n_0;
    wire memAWrite[11]_i_10_n_0;
    wire memAWrite[11]_i_11_n_0;
    wire memAWrite[11]_i_12_n_0;
    wire memAWrite[11]_i_2_n_0;
    wire memAWrite[11]_i_3_n_0;
    wire memAWrite[11]_i_5_n_0;
    wire memAWrite[11]_i_6_n_0;
    wire memAWrite[11]_i_9_n_0;
    wire memAWrite[12]_i_2_n_0;
    wire memAWrite[12]_i_3_n_0;
    wire memAWrite[12]_i_5_n_0;
    wire memAWrite[12]_i_6_n_0;
    wire memAWrite[13]_i_2_n_0;
    wire memAWrite[13]_i_3_n_0;
    wire memAWrite[13]_i_5_n_0;
    wire memAWrite[13]_i_6_n_0;
    wire memAWrite[14]_i_2_n_0;
    wire memAWrite[14]_i_3_n_0;
    wire memAWrite[14]_i_5_n_0;
    wire memAWrite[14]_i_6_n_0;
    wire memAWrite[15]_i_2_n_0;
    wire memAWrite[15]_i_3_n_0;
    wire memAWrite[15]_i_4_n_0;
    wire memAWrite[15]_i_6_n_0;
    wire memAWrite[15]_i_7_n_0;
    wire memAWrite[15]_i_8_n_0;
    wire memAWrite[15]_i_9_n_0;
    wire memAWrite[16]_i_2_n_0;
    wire memAWrite[16]_i_3_n_0;
    wire memAWrite[16]_i_4_n_0;
    wire memAWrite[17]_i_2_n_0;
    wire memAWrite[17]_i_3_n_0;
    wire memAWrite[17]_i_4_n_0;
    wire memAWrite[18]_i_2_n_0;
    wire memAWrite[18]_i_3_n_0;
    wire memAWrite[18]_i_4_n_0;
    wire memAWrite[19]_i_2_n_0;
    wire memAWrite[19]_i_3_n_0;
    wire memAWrite[19]_i_4_n_0;
    wire memAWrite[19]_i_6_n_0;
    wire memAWrite[19]_i_7_n_0;
    wire memAWrite[19]_i_8_n_0;
    wire memAWrite[19]_i_9_n_0;
    wire memAWrite[1]_i_2_n_0;
    wire memAWrite[1]_i_3_n_0;
    wire memAWrite[1]_i_5_n_0;
    wire memAWrite[20]_i_2_n_0;
    wire memAWrite[20]_i_3_n_0;
    wire memAWrite[20]_i_4_n_0;
    wire memAWrite[21]_i_2_n_0;
    wire memAWrite[21]_i_3_n_0;
    wire memAWrite[21]_i_4_n_0;
    wire memAWrite[22]_i_2_n_0;
    wire memAWrite[22]_i_3_n_0;
    wire memAWrite[22]_i_4_n_0;
    wire memAWrite[23]_i_2_n_0;
    wire memAWrite[23]_i_3_n_0;
    wire memAWrite[23]_i_4_n_0;
    wire memAWrite[23]_i_6_n_0;
    wire memAWrite[23]_i_7_n_0;
    wire memAWrite[23]_i_8_n_0;
    wire memAWrite[23]_i_9_n_0;
    wire memAWrite[24]_i_2_n_0;
    wire memAWrite[24]_i_3_n_0;
    wire memAWrite[24]_i_4_n_0;
    wire memAWrite[25]_i_2_n_0;
    wire memAWrite[25]_i_3_n_0;
    wire memAWrite[25]_i_4_n_0;
    wire memAWrite[26]_i_2_n_0;
    wire memAWrite[26]_i_3_n_0;
    wire memAWrite[26]_i_4_n_0;
    wire memAWrite[27]_i_2_n_0;
    wire memAWrite[27]_i_3_n_0;
    wire memAWrite[27]_i_4_n_0;
    wire memAWrite[27]_i_6_n_0;
    wire memAWrite[27]_i_7_n_0;
    wire memAWrite[27]_i_8_n_0;
    wire memAWrite[27]_i_9_n_0;
    wire memAWrite[28]_i_2_n_0;
    wire memAWrite[28]_i_3_n_0;
    wire memAWrite[28]_i_4_n_0;
    wire memAWrite[29]_i_2_n_0;
    wire memAWrite[29]_i_3_n_0;
    wire memAWrite[29]_i_4_n_0;
    wire memAWrite[2]_i_2_n_0;
    wire memAWrite[2]_i_3_n_0;
    wire memAWrite[2]_i_6_n_0;
    wire memAWrite[30]_i_2_n_0;
    wire memAWrite[30]_i_3_n_0;
    wire memAWrite[30]_i_4_n_0;
    wire memAWrite[31]_i_10_n_0;
    wire memAWrite[31]_i_2_n_0;
    wire memAWrite[31]_i_3_n_0;
    wire memAWrite[31]_i_5_n_0;
    wire memAWrite[31]_i_7_n_0;
    wire memAWrite[31]_i_8_n_0;
    wire memAWrite[31]_i_9_n_0;
    wire memAWrite[3]_i_10_n_0;
    wire memAWrite[3]_i_11_n_0;
    wire memAWrite[3]_i_2_n_0;
    wire memAWrite[3]_i_3_n_0;
    wire memAWrite[3]_i_6_n_0;
    wire memAWrite[3]_i_8_n_0;
    wire memAWrite[3]_i_9_n_0;
    wire memAWrite[4]_i_2_n_0;
    wire memAWrite[4]_i_3_n_0;
    wire memAWrite[4]_i_6_n_0;
    wire memAWrite[5]_i_2_n_0;
    wire memAWrite[5]_i_3_n_0;
    wire memAWrite[5]_i_6_n_0;
    wire memAWrite[6]_i_2_n_0;
    wire memAWrite[6]_i_3_n_0;
    wire memAWrite[6]_i_6_n_0;
    wire memAWrite[7]_i_10_n_0;
    wire memAWrite[7]_i_11_n_0;
    wire memAWrite[7]_i_12_n_0;
    wire memAWrite[7]_i_2_n_0;
    wire memAWrite[7]_i_3_n_0;
    wire memAWrite[7]_i_5_n_0;
    wire memAWrite[7]_i_6_n_0;
    wire memAWrite[7]_i_9_n_0;
    wire memAWrite[8]_i_2_n_0;
    wire memAWrite[8]_i_3_n_0;
    wire memAWrite[8]_i_5_n_0;
    wire memAWrite[8]_i_6_n_0;
    wire memAWrite[9]_i_2_n_0;
    wire memAWrite[9]_i_3_n_0;
    wire memAWrite[9]_i_5_n_0;
    wire memAWrite[9]_i_6_n_0;
    wire memAWrite_reg[11]_i_8_n_0;
    wire memAWrite_reg[11]_i_8_n_1;
    wire memAWrite_reg[11]_i_8_n_2;
    wire memAWrite_reg[11]_i_8_n_3;
    wire memAWrite_reg[11]_i_8_n_4;
    wire memAWrite_reg[11]_i_8_n_5;
    wire memAWrite_reg[11]_i_8_n_6;
    wire memAWrite_reg[11]_i_8_n_7;
    wire memAWrite_reg[15]_i_5_n_0;
    wire memAWrite_reg[15]_i_5_n_1;
    wire memAWrite_reg[15]_i_5_n_2;
    wire memAWrite_reg[15]_i_5_n_3;
    wire memAWrite_reg[15]_i_5_n_4;
    wire memAWrite_reg[15]_i_5_n_5;
    wire memAWrite_reg[15]_i_5_n_6;
    wire memAWrite_reg[15]_i_5_n_7;
    wire memAWrite_reg[19]_i_5_n_0;
    wire memAWrite_reg[19]_i_5_n_1;
    wire memAWrite_reg[19]_i_5_n_2;
    wire memAWrite_reg[19]_i_5_n_3;
    wire memAWrite_reg[19]_i_5_n_4;
    wire memAWrite_reg[19]_i_5_n_5;
    wire memAWrite_reg[19]_i_5_n_6;
    wire memAWrite_reg[19]_i_5_n_7;
    wire memAWrite_reg[23]_i_5_n_0;
    wire memAWrite_reg[23]_i_5_n_1;
    wire memAWrite_reg[23]_i_5_n_2;
    wire memAWrite_reg[23]_i_5_n_3;
    wire memAWrite_reg[23]_i_5_n_4;
    wire memAWrite_reg[23]_i_5_n_5;
    wire memAWrite_reg[23]_i_5_n_6;
    wire memAWrite_reg[23]_i_5_n_7;
    wire memAWrite_reg[27]_i_5_n_0;
    wire memAWrite_reg[27]_i_5_n_1;
    wire memAWrite_reg[27]_i_5_n_2;
    wire memAWrite_reg[27]_i_5_n_3;
    wire memAWrite_reg[27]_i_5_n_4;
    wire memAWrite_reg[27]_i_5_n_5;
    wire memAWrite_reg[27]_i_5_n_6;
    wire memAWrite_reg[27]_i_5_n_7;
    wire [31:0]memAWrite_reg[31];
    wire [31:0]memAWrite_reg[31]_0;
    wire memAWrite_reg[31]_i_6_n_1;
    wire memAWrite_reg[31]_i_6_n_2;
    wire memAWrite_reg[31]_i_6_n_3;
    wire memAWrite_reg[31]_i_6_n_4;
    wire memAWrite_reg[31]_i_6_n_5;
    wire memAWrite_reg[31]_i_6_n_6;
    wire memAWrite_reg[31]_i_6_n_7;
    wire memAWrite_reg[3]_i_7_n_0;
    wire memAWrite_reg[3]_i_7_n_1;
    wire memAWrite_reg[3]_i_7_n_2;
    wire memAWrite_reg[3]_i_7_n_3;
    wire memAWrite_reg[3]_i_7_n_4;
    wire memAWrite_reg[3]_i_7_n_5;
    wire memAWrite_reg[3]_i_7_n_6;
    wire memAWrite_reg[3]_i_7_n_7;
    wire memAWrite_reg[7]_i_8_n_0;
    wire memAWrite_reg[7]_i_8_n_1;
    wire memAWrite_reg[7]_i_8_n_2;
    wire memAWrite_reg[7]_i_8_n_3;
    wire memAWrite_reg[7]_i_8_n_4;
    wire memAWrite_reg[7]_i_8_n_5;
    wire memAWrite_reg[7]_i_8_n_6;
    wire memAWrite_reg[7]_i_8_n_7;
    wire [12:0]memBAddr_reg[14];
    wire [31:0]memBRead;
    wire memBWriteEnable;
    wire [31:0]memBWrite_reg[31];
    wire [31:0]mem_read_IBUF;
    wire [6:0]opcode_reg;
    wire opcode_reg[0]_0;
    wire opcode_reg[0]_1;
    wire opcode_reg[1]_0;
    wire [4:0]opcode_reg[6]_0;
    wire [3:0]out;
    wire out_mem_readEnable_reg;
    wire [13:2]pc_reg;
    wire [14:0]pc_reg[14];
    wire pc_reg[14]_0;
    wire [13:0]pc_reg[14]_1;
    wire [1:0]pc_reg[1];
    wire sp[10]_i_2_n_0;
    wire sp[11]_i_2_n_0;
    wire sp[12]_i_2_n_0;
    wire sp[13]_i_2_n_0;
    wire sp[14]_i_3_n_0;
    wire sp[2]_i_3_n_0;
    wire sp[3]_i_2_n_0;
    wire sp[4]_i_2_n_0;
    wire sp[5]_i_2_n_0;
    wire sp[6]_i_2_n_0;
    wire sp[7]_i_2_n_0;
    wire sp[8]_i_2_n_0;
    wire sp[9]_i_2_n_0;
    wire [3:0]sp_reg[10];
    wire [12:0]sp_reg[14];
    wire [12:0]sp_reg[14]_0;
    wire [3:0]sp_reg[2];

    LUT6 FSM_sequential_state[1]_i_1
    (
        .O(D[0]),
        .I0(in_mem_busy_IBUF),
        .I1(FSM_sequential_state[1]_i_2_n_0),
        .I2(out[2]),
        .I3(out[1]),
        .I4(out[0]),
        .I5(out[3])
    );
    LUT5 FSM_sequential_state[1]_i_2
    (
        .O(FSM_sequential_state[1]_i_2_n_0),
        .I0(out[0]),
        .I1(FSM_sequential_state_reg[2]),
        .I2(Q[3]),
        .I3(memARead[15]),
        .I4(Q[1])
    );
    LUT5 FSM_sequential_state[2]_i_1
    (
        .O(D[1]),
        .I0(FSM_sequential_state[2]_i_2_n_0),
        .I1(FSM_sequential_state_reg[0]),
        .I2(out[1]),
        .I3(out[2]),
        .I4(out[3])
    );
    LUT6 FSM_sequential_state[2]_i_2
    (
        .O(FSM_sequential_state[2]_i_2_n_0),
        .I0(out[0]),
        .I1(Q[3]),
        .I2(Q[0]),
        .I3(Q[2]),
        .I4(memARead[15]),
        .I5(Q[1])
    );
    LUT6 FSM_sequential_state[3]_i_2
    (
        .O(D[2]),
        .I0(FSM_sequential_state_reg[3]),
        .I1(FSM_sequential_state[3]_i_4_n_0),
        .I2(Q[2]),
        .I3(Q[4]),
        .I4(Q[3]),
        .I5(FSM_sequential_state_reg[1])
    );
    LUT4 FSM_sequential_state[3]_i_4
    (
        .O(FSM_sequential_state[3]_i_4_n_0),
        .I0(Q[1]),
        .I1(Q[2]),
        .I2(memARead[15]),
        .I3(Q[0])
    );
    GND GND
    (
        .G(<const0>)
    );
    VCC VCC
    (
        .P(<const1>)
    );
    LUT6 decodedOpcode[0]_i_1
    (
        .O(decodedOpcode_reg[4][0]),
        .I0(FSM_sequential_state_reg[1]_0),
        .I1(decodedOpcode[4]_i_4_n_0),
        .I2(opcode_reg[6]),
        .I3(opcode_reg[5]),
        .I4(decodedOpcode[0]_i_2_n_0),
        .I5(inInterrupt_reg)
    );
    LUT5 decodedOpcode[0]_i_2
    (
        .O(decodedOpcode[0]_i_2_n_0),
        .I0(opcode_reg[4]),
        .I1(opcode_reg[2]),
        .I2(opcode_reg[0]),
        .I3(opcode_reg[3]),
        .I4(opcode_reg[1])
    );
    LUT6 decodedOpcode[1]_i_1
    (
        .O(decodedOpcode_reg[4][1]),
        .I0(FSM_sequential_state_reg[1]_0),
        .I1(decodedOpcode[1]_i_2_n_0),
        .I2(decodedOpcode[3]_i_2_n_0),
        .I3(opcode_reg[5]),
        .I4(decodedOpcode[4]_i_4_n_0),
        .I5(inInterrupt_reg)
    );
    LUT5 decodedOpcode[1]_i_2
    (
        .O(decodedOpcode[1]_i_2_n_0),
        .I0(opcode_reg[5]),
        .I1(opcode_reg[2]),
        .I2(opcode_reg[3]),
        .I3(opcode_reg[1]),
        .I4(opcode_reg[0])
    );
    LUT5 decodedOpcode[2]_i_1
    (
        .O(decodedOpcode_reg[4][2]),
        .I0(FSM_sequential_state_reg[1]_0),
        .I1(inInterrupt_reg),
        .I2(decodedOpcode[2]_i_2_n_0),
        .I3(decodedOpcode[2]_i_3_n_0),
        .I4(decodedOpcode[2]_i_4_n_0)
    );
    LUT3 decodedOpcode[2]_i_2
    (
        .O(decodedOpcode[2]_i_2_n_0),
        .I0(decodedOpcode[4]_i_4_n_0),
        .I1(opcode_reg[6]),
        .I2(opcode_reg[5])
    );
    LUT4 decodedOpcode[2]_i_3
    (
        .O(decodedOpcode[2]_i_3_n_0),
        .I0(opcode_reg[3]),
        .I1(opcode_reg[0]),
        .I2(opcode_reg[1]),
        .I3(opcode_reg[2])
    );
    LUT6 decodedOpcode[2]_i_4
    (
        .O(decodedOpcode[2]_i_4_n_0),
        .I0(opcode_reg[4]),
        .I1(opcode_reg[1]),
        .I2(opcode_reg[3]),
        .I3(opcode_reg[2]),
        .I4(opcode_reg[6]),
        .I5(opcode_reg[5])
    );
    LUT5 decodedOpcode[3]_i_1
    (
        .O(decodedOpcode_reg[4][3]),
        .I0(FSM_sequential_state_reg[1]_0),
        .I1(opcode_reg[5]),
        .I2(decodedOpcode[3]_i_2_n_0),
        .I3(decodedOpcode[3]_i_3_n_0),
        .I4(inInterrupt_reg)
    );
    LUT2 decodedOpcode[3]_i_2
    (
        .O(decodedOpcode[3]_i_2_n_0),
        .I0(opcode_reg[4]),
        .I1(opcode_reg[6])
    );
    LUT5 decodedOpcode[3]_i_3
    (
        .O(decodedOpcode[3]_i_3_n_0),
        .I0(opcode_reg[0]),
        .I1(opcode_reg[1]),
        .I2(opcode_reg[2]),
        .I3(opcode_reg[3]),
        .I4(decodedOpcode[4]_i_4_n_0)
    );
    LUT5 decodedOpcode[4]_i_1
    (
        .O(decodedOpcode_reg[4][4]),
        .I0(FSM_sequential_state_reg[1]_0),
        .I1(decodedOpcode[4]_i_3_n_0),
        .I2(decodedOpcode[4]_i_4_n_0),
        .I3(opcode_reg[5]),
        .I4(inInterrupt_reg)
    );
    LUT5 decodedOpcode[4]_i_3
    (
        .O(decodedOpcode[4]_i_3_n_0),
        .I0(opcode_reg[4]),
        .I1(opcode_reg[6]),
        .I2(opcode_reg[3]),
        .I3(opcode_reg[1]),
        .I4(opcode_reg[2])
    );
    LUT6 decodedOpcode[4]_i_4
    (
        .O(decodedOpcode[4]_i_4_n_0),
        .I0(memBRead[15]),
        .I1(memBRead[7]),
        .I2(pc_reg[1][1]),
        .I3(pc_reg[1][0]),
        .I4(memBRead[31]),
        .I5(memBRead[23])
    );
    LUT6 memAAddr[10]_i_1
    (
        .O(memAAddr_reg[14][8]),
        .I0(memARead[10]),
        .I1(out[3]),
        .I2(out[1]),
        .I3(out[2]),
        .I4(memAAddr[10]_i_2_n_0),
        .I5(sp_reg[14]_0[8])
    );
    LUT6 memAAddr[10]_i_2
    (
        .O(memAAddr[10]_i_2_n_0),
        .I0(memAAddr[10]_i_3_n_0),
        .I1(decodedOpcode_reg[4]_1),
        .I2(sp_reg[14]_0[8]),
        .I3(decodedOpcode_reg[1]),
        .I4(sp_reg[10][3]),
        .I5(decodedOpcode_reg[2]_13)
    );
    LUT5 memAAddr[10]_i_3
    (
        .O(memAAddr[10]_i_3_n_0),
        .I0(Q[1]),
        .I1(Q[2]),
        .I2(Q[3]),
        .I3(Q[0]),
        .I4(memARead[10])
    );
    LUT6 memAAddr[11]_i_1
    (
        .O(memAAddr_reg[14][9]),
        .I0(memARead[11]),
        .I1(out[3]),
        .I2(out[1]),
        .I3(out[2]),
        .I4(memAAddr[11]_i_2_n_0),
        .I5(sp_reg[14]_0[9])
    );
    LUT6 memAAddr[11]_i_2
    (
        .O(memAAddr[11]_i_2_n_0),
        .I0(memAAddr[11]_i_3_n_0),
        .I1(decodedOpcode_reg[4]_1),
        .I2(sp_reg[14]_0[9]),
        .I3(decodedOpcode_reg[1]),
        .I4(O[0]),
        .I5(decodedOpcode_reg[2]_14)
    );
    LUT5 memAAddr[11]_i_3
    (
        .O(memAAddr[11]_i_3_n_0),
        .I0(Q[1]),
        .I1(Q[2]),
        .I2(Q[3]),
        .I3(Q[0]),
        .I4(memARead[11])
    );
    LUT6 memAAddr[12]_i_1
    (
        .O(memAAddr_reg[14][10]),
        .I0(memARead[12]),
        .I1(out[3]),
        .I2(out[1]),
        .I3(out[2]),
        .I4(memAAddr[12]_i_2_n_0),
        .I5(sp_reg[14]_0[10])
    );
    LUT6 memAAddr[12]_i_2
    (
        .O(memAAddr[12]_i_2_n_0),
        .I0(memAAddr[12]_i_3_n_0),
        .I1(decodedOpcode_reg[4]_1),
        .I2(sp_reg[14]_0[10]),
        .I3(decodedOpcode_reg[1]),
        .I4(O[1]),
        .I5(decodedOpcode_reg[2]_15)
    );
    LUT5 memAAddr[12]_i_3
    (
        .O(memAAddr[12]_i_3_n_0),
        .I0(Q[1]),
        .I1(Q[2]),
        .I2(Q[3]),
        .I3(Q[0]),
        .I4(memARead[12])
    );
    LUT6 memAAddr[13]_i_1
    (
        .O(memAAddr_reg[14][11]),
        .I0(memARead[13]),
        .I1(out[3]),
        .I2(out[1]),
        .I3(out[2]),
        .I4(memAAddr[13]_i_2_n_0),
        .I5(sp_reg[14]_0[11])
    );
    LUT6 memAAddr[13]_i_2
    (
        .O(memAAddr[13]_i_2_n_0),
        .I0(memAAddr[13]_i_3_n_0),
        .I1(decodedOpcode_reg[4]_1),
        .I2(sp_reg[14]_0[11]),
        .I3(decodedOpcode_reg[1]),
        .I4(O[2]),
        .I5(decodedOpcode_reg[2]_16)
    );
    LUT5 memAAddr[13]_i_3
    (
        .O(memAAddr[13]_i_3_n_0),
        .I0(Q[1]),
        .I1(Q[2]),
        .I2(Q[3]),
        .I3(Q[0]),
        .I4(memARead[13])
    );
    LUT6 memAAddr[14]_i_1
    (
        .O(memAAddr_reg[14][12]),
        .I0(memARead[14]),
        .I1(out[3]),
        .I2(out[1]),
        .I3(out[2]),
        .I4(memAAddr[14]_i_2_n_0),
        .I5(sp_reg[14]_0[12])
    );
    LUT6 memAAddr[14]_i_2
    (
        .O(memAAddr[14]_i_2_n_0),
        .I0(memAAddr[14]_i_3_n_0),
        .I1(decodedOpcode_reg[4]_1),
        .I2(sp_reg[14]_0[12]),
        .I3(decodedOpcode_reg[1]),
        .I4(O[3]),
        .I5(decodedOpcode_reg[2]_17)
    );
    LUT5 memAAddr[14]_i_3
    (
        .O(memAAddr[14]_i_3_n_0),
        .I0(Q[1]),
        .I1(Q[2]),
        .I2(Q[3]),
        .I3(Q[0]),
        .I4(memARead[14])
    );
    LUT6 memAAddr[2]_i_1
    (
        .O(memAAddr_reg[14][0]),
        .I0(memARead[2]),
        .I1(out[3]),
        .I2(out[1]),
        .I3(out[2]),
        .I4(memAAddr[2]_i_2_n_0),
        .I5(sp_reg[14]_0[0])
    );
    LUT6 memAAddr[2]_i_2
    (
        .O(memAAddr[2]_i_2_n_0),
        .I0(decodedOpcode_reg[0]_3),
        .I1(memARead[2]),
        .I2(decodedOpcode_reg[4]_1),
        .I3(decodedOpcode_reg[1]),
        .I4(sp_reg[14]_0[0]),
        .I5(decodedOpcode_reg[2]_5)
    );
    LUT6 memAAddr[3]_i_1
    (
        .O(memAAddr_reg[14][1]),
        .I0(memARead[3]),
        .I1(out[3]),
        .I2(out[1]),
        .I3(out[2]),
        .I4(memAAddr[3]_i_2_n_0),
        .I5(sp_reg[14]_0[1])
    );
    LUT6 memAAddr[3]_i_2
    (
        .O(memAAddr[3]_i_2_n_0),
        .I0(memAAddr[3]_i_3_n_0),
        .I1(decodedOpcode_reg[4]_1),
        .I2(sp_reg[14]_0[1]),
        .I3(decodedOpcode_reg[1]),
        .I4(sp_reg[2][0]),
        .I5(decodedOpcode_reg[2]_6)
    );
    LUT5 memAAddr[3]_i_3
    (
        .O(memAAddr[3]_i_3_n_0),
        .I0(Q[1]),
        .I1(Q[2]),
        .I2(Q[3]),
        .I3(Q[0]),
        .I4(memARead[3])
    );
    LUT6 memAAddr[4]_i_1
    (
        .O(memAAddr_reg[14][2]),
        .I0(memARead[4]),
        .I1(out[3]),
        .I2(out[1]),
        .I3(out[2]),
        .I4(memAAddr[4]_i_2_n_0),
        .I5(sp_reg[14]_0[2])
    );
    LUT6 memAAddr[4]_i_2
    (
        .O(memAAddr[4]_i_2_n_0),
        .I0(memAAddr[4]_i_3_n_0),
        .I1(decodedOpcode_reg[4]_1),
        .I2(sp_reg[14]_0[2]),
        .I3(decodedOpcode_reg[1]),
        .I4(sp_reg[2][1]),
        .I5(decodedOpcode_reg[2]_7)
    );
    LUT5 memAAddr[4]_i_3
    (
        .O(memAAddr[4]_i_3_n_0),
        .I0(Q[1]),
        .I1(Q[2]),
        .I2(Q[3]),
        .I3(Q[0]),
        .I4(memARead[4])
    );
    LUT6 memAAddr[5]_i_1
    (
        .O(memAAddr_reg[14][3]),
        .I0(memARead[5]),
        .I1(out[3]),
        .I2(out[1]),
        .I3(out[2]),
        .I4(memAAddr[5]_i_2_n_0),
        .I5(sp_reg[14]_0[3])
    );
    LUT6 memAAddr[5]_i_2
    (
        .O(memAAddr[5]_i_2_n_0),
        .I0(memAAddr[5]_i_3_n_0),
        .I1(decodedOpcode_reg[4]_1),
        .I2(sp_reg[14]_0[3]),
        .I3(decodedOpcode_reg[1]),
        .I4(sp_reg[2][2]),
        .I5(decodedOpcode_reg[2]_8)
    );
    LUT5 memAAddr[5]_i_3
    (
        .O(memAAddr[5]_i_3_n_0),
        .I0(Q[1]),
        .I1(Q[2]),
        .I2(Q[3]),
        .I3(Q[0]),
        .I4(memARead[5])
    );
    LUT6 memAAddr[6]_i_1
    (
        .O(memAAddr_reg[14][4]),
        .I0(memARead[6]),
        .I1(out[3]),
        .I2(out[1]),
        .I3(out[2]),
        .I4(memAAddr[6]_i_2_n_0),
        .I5(sp_reg[14]_0[4])
    );
    LUT6 memAAddr[6]_i_2
    (
        .O(memAAddr[6]_i_2_n_0),
        .I0(memAAddr[6]_i_3_n_0),
        .I1(decodedOpcode_reg[4]_1),
        .I2(sp_reg[14]_0[4]),
        .I3(decodedOpcode_reg[1]),
        .I4(sp_reg[2][3]),
        .I5(decodedOpcode_reg[2]_9)
    );
    LUT5 memAAddr[6]_i_3
    (
        .O(memAAddr[6]_i_3_n_0),
        .I0(Q[1]),
        .I1(Q[2]),
        .I2(Q[3]),
        .I3(Q[0]),
        .I4(memARead[6])
    );
    LUT6 memAAddr[7]_i_1
    (
        .O(memAAddr_reg[14][5]),
        .I0(memARead[7]),
        .I1(out[3]),
        .I2(out[1]),
        .I3(out[2]),
        .I4(memAAddr[7]_i_2_n_0),
        .I5(sp_reg[14]_0[5])
    );
    LUT6 memAAddr[7]_i_2
    (
        .O(memAAddr[7]_i_2_n_0),
        .I0(memAAddr[7]_i_3_n_0),
        .I1(decodedOpcode_reg[4]_1),
        .I2(sp_reg[14]_0[5]),
        .I3(decodedOpcode_reg[1]),
        .I4(sp_reg[10][0]),
        .I5(decodedOpcode_reg[2]_10)
    );
    LUT5 memAAddr[7]_i_3
    (
        .O(memAAddr[7]_i_3_n_0),
        .I0(Q[1]),
        .I1(Q[2]),
        .I2(Q[3]),
        .I3(Q[0]),
        .I4(memARead[7])
    );
    LUT6 memAAddr[8]_i_1
    (
        .O(memAAddr_reg[14][6]),
        .I0(memARead[8]),
        .I1(out[3]),
        .I2(out[1]),
        .I3(out[2]),
        .I4(memAAddr[8]_i_2_n_0),
        .I5(sp_reg[14]_0[6])
    );
    LUT6 memAAddr[8]_i_2
    (
        .O(memAAddr[8]_i_2_n_0),
        .I0(memAAddr[8]_i_3_n_0),
        .I1(decodedOpcode_reg[4]_1),
        .I2(sp_reg[14]_0[6]),
        .I3(decodedOpcode_reg[1]),
        .I4(sp_reg[10][1]),
        .I5(decodedOpcode_reg[2]_11)
    );
    LUT5 memAAddr[8]_i_3
    (
        .O(memAAddr[8]_i_3_n_0),
        .I0(Q[1]),
        .I1(Q[2]),
        .I2(Q[3]),
        .I3(Q[0]),
        .I4(memARead[8])
    );
    LUT6 memAAddr[9]_i_1
    (
        .O(memAAddr_reg[14][7]),
        .I0(memARead[9]),
        .I1(out[3]),
        .I2(out[1]),
        .I3(out[2]),
        .I4(memAAddr[9]_i_2_n_0),
        .I5(sp_reg[14]_0[7])
    );
    LUT6 memAAddr[9]_i_2
    (
        .O(memAAddr[9]_i_2_n_0),
        .I0(memAAddr[9]_i_3_n_0),
        .I1(decodedOpcode_reg[4]_1),
        .I2(sp_reg[14]_0[7]),
        .I3(decodedOpcode_reg[1]),
        .I4(sp_reg[10][2]),
        .I5(decodedOpcode_reg[2]_12)
    );
    LUT5 memAAddr[9]_i_3
    (
        .O(memAAddr[9]_i_3_n_0),
        .I0(Q[1]),
        .I1(Q[2]),
        .I2(Q[3]),
        .I3(Q[0]),
        .I4(memARead[9])
    );
    LUT6 memAWrite[0]_i_1
    (
        .O(memAWrite_reg[31][0]),
        .I0(memBRead[0]),
        .I1(out[3]),
        .I2(memAWrite[0]_i_2_n_0),
        .I3(out[1]),
        .I4(out[2]),
        .I5(memAWrite[0]_i_3_n_0)
    );
    LUT6 memAWrite[0]_i_2
    (
        .O(memAWrite[0]_i_2_n_0),
        .I0(memARead[0]),
        .I1(out[1]),
        .I2(decodedOpcode_reg[2]),
        .I3(memARead[31]),
        .I4(opcode_reg[0]_0),
        .I5(memAWrite[0]_i_5_n_0)
    );
    LUT6 memAWrite[0]_i_3
    (
        .O(memAWrite[0]_i_3_n_0),
        .I0(mem_read_IBUF[0]),
        .I1(out[0]),
        .I2(memAWrite_reg[3]_i_7_n_7),
        .I3(out[1]),
        .I4(memBRead[0]),
        .I5(memARead[0])
    );
    LUT5 memAWrite[0]_i_5
    (
        .O(memAWrite[0]_i_5_n_0),
        .I0(memARead[0]),
        .I1(Q[0]),
        .I2(pc_reg[1][0]),
        .I3(Q[2]),
        .I4(Q[3])
    );
    LUT6 memAWrite[10]_i_1
    (
        .O(memAWrite_reg[31][10]),
        .I0(memBRead[10]),
        .I1(out[3]),
        .I2(memAWrite[10]_i_2_n_0),
        .I3(out[1]),
        .I4(out[2]),
        .I5(memAWrite[10]_i_3_n_0)
    );
    LUT6 memAWrite[10]_i_2
    (
        .O(memAWrite[10]_i_2_n_0),
        .I0(memARead[10]),
        .I1(out[1]),
        .I2(pc_reg[10]),
        .I3(memAWrite[10]_i_5_n_0),
        .I4(memAWrite[10]_i_6_n_0),
        .I5(decodedOpcode_reg[3]_3)
    );
    LUT6 memAWrite[10]_i_3
    (
        .O(memAWrite[10]_i_3_n_0),
        .I0(mem_read_IBUF[10]),
        .I1(out[0]),
        .I2(memAWrite_reg[11]_i_8_n_5),
        .I3(out[1]),
        .I4(memBRead[10]),
        .I5(memARead[10])
    );
    LUT6 memAWrite[10]_i_5
    (
        .O(memAWrite[10]_i_5_n_0),
        .I0(memARead[10]),
        .I1(Q[3]),
        .I2(memARead[3]),
        .I3(Q[2]),
        .I4(Q[0]),
        .I5(idim_flag)
    );
    LUT4 memAWrite[10]_i_6
    (
        .O(memAWrite[10]_i_6_n_0),
        .I0(Q[0]),
        .I1(Q[3]),
        .I2(Q[2]),
        .I3(memARead[21])
    );
    LUT6 memAWrite[11]_i_1
    (
        .O(memAWrite_reg[31][11]),
        .I0(memBRead[11]),
        .I1(out[3]),
        .I2(memAWrite[11]_i_2_n_0),
        .I3(out[1]),
        .I4(out[2]),
        .I5(memAWrite[11]_i_3_n_0)
    );
    LUT2 memAWrite[11]_i_10
    (
        .O(memAWrite[11]_i_10_n_0),
        .I0(memARead[10]),
        .I1(memBRead[10])
    );
    LUT2 memAWrite[11]_i_11
    (
        .O(memAWrite[11]_i_11_n_0),
        .I0(memARead[9]),
        .I1(memBRead[9])
    );
    LUT2 memAWrite[11]_i_12
    (
        .O(memAWrite[11]_i_12_n_0),
        .I0(memARead[8]),
        .I1(memBRead[8])
    );
    LUT6 memAWrite[11]_i_2
    (
        .O(memAWrite[11]_i_2_n_0),
        .I0(memARead[11]),
        .I1(out[1]),
        .I2(pc_reg[11]),
        .I3(memAWrite[11]_i_5_n_0),
        .I4(memAWrite[11]_i_6_n_0),
        .I5(decodedOpcode_reg[3]_2)
    );
    LUT6 memAWrite[11]_i_3
    (
        .O(memAWrite[11]_i_3_n_0),
        .I0(mem_read_IBUF[11]),
        .I1(out[0]),
        .I2(memAWrite_reg[11]_i_8_n_4),
        .I3(out[1]),
        .I4(memBRead[11]),
        .I5(memARead[11])
    );
    LUT6 memAWrite[11]_i_5
    (
        .O(memAWrite[11]_i_5_n_0),
        .I0(memARead[11]),
        .I1(Q[3]),
        .I2(memARead[4]),
        .I3(Q[2]),
        .I4(Q[0]),
        .I5(idim_flag)
    );
    LUT4 memAWrite[11]_i_6
    (
        .O(memAWrite[11]_i_6_n_0),
        .I0(Q[0]),
        .I1(Q[3]),
        .I2(Q[2]),
        .I3(memARead[20])
    );
    LUT2 memAWrite[11]_i_9
    (
        .O(memAWrite[11]_i_9_n_0),
        .I0(memARead[11]),
        .I1(memBRead[11])
    );
    LUT6 memAWrite[12]_i_1
    (
        .O(memAWrite_reg[31][12]),
        .I0(memBRead[12]),
        .I1(out[3]),
        .I2(memAWrite[12]_i_2_n_0),
        .I3(out[1]),
        .I4(out[2]),
        .I5(memAWrite[12]_i_3_n_0)
    );
    LUT6 memAWrite[12]_i_2
    (
        .O(memAWrite[12]_i_2_n_0),
        .I0(memARead[12]),
        .I1(out[1]),
        .I2(pc_reg[12]),
        .I3(memAWrite[12]_i_5_n_0),
        .I4(memAWrite[12]_i_6_n_0),
        .I5(decodedOpcode_reg[3]_1)
    );
    LUT6 memAWrite[12]_i_3
    (
        .O(memAWrite[12]_i_3_n_0),
        .I0(mem_read_IBUF[12]),
        .I1(out[0]),
        .I2(memAWrite_reg[15]_i_5_n_7),
        .I3(out[1]),
        .I4(memBRead[12]),
        .I5(memARead[12])
    );
    LUT6 memAWrite[12]_i_5
    (
        .O(memAWrite[12]_i_5_n_0),
        .I0(memARead[12]),
        .I1(Q[3]),
        .I2(memARead[5]),
        .I3(Q[2]),
        .I4(Q[0]),
        .I5(idim_flag)
    );
    LUT4 memAWrite[12]_i_6
    (
        .O(memAWrite[12]_i_6_n_0),
        .I0(Q[0]),
        .I1(Q[3]),
        .I2(Q[2]),
        .I3(memARead[19])
    );
    LUT6 memAWrite[13]_i_1
    (
        .O(memAWrite_reg[31][13]),
        .I0(memBRead[13]),
        .I1(out[3]),
        .I2(memAWrite[13]_i_2_n_0),
        .I3(out[1]),
        .I4(out[2]),
        .I5(memAWrite[13]_i_3_n_0)
    );
    LUT6 memAWrite[13]_i_2
    (
        .O(memAWrite[13]_i_2_n_0),
        .I0(memARead[13]),
        .I1(out[1]),
        .I2(pc_reg[13]),
        .I3(memAWrite[13]_i_5_n_0),
        .I4(memAWrite[13]_i_6_n_0),
        .I5(decodedOpcode_reg[3]_0)
    );
    LUT6 memAWrite[13]_i_3
    (
        .O(memAWrite[13]_i_3_n_0),
        .I0(mem_read_IBUF[13]),
        .I1(out[0]),
        .I2(memAWrite_reg[15]_i_5_n_6),
        .I3(out[1]),
        .I4(memBRead[13]),
        .I5(memARead[13])
    );
    LUT6 memAWrite[13]_i_5
    (
        .O(memAWrite[13]_i_5_n_0),
        .I0(memARead[13]),
        .I1(Q[3]),
        .I2(memARead[6]),
        .I3(Q[2]),
        .I4(Q[0]),
        .I5(idim_flag)
    );
    LUT4 memAWrite[13]_i_6
    (
        .O(memAWrite[13]_i_6_n_0),
        .I0(Q[0]),
        .I1(Q[3]),
        .I2(Q[2]),
        .I3(memARead[18])
    );
    LUT6 memAWrite[14]_i_1
    (
        .O(memAWrite_reg[31][14]),
        .I0(memBRead[14]),
        .I1(out[3]),
        .I2(memAWrite[14]_i_2_n_0),
        .I3(out[1]),
        .I4(out[2]),
        .I5(memAWrite[14]_i_3_n_0)
    );
    LUT6 memAWrite[14]_i_2
    (
        .O(memAWrite[14]_i_2_n_0),
        .I0(memARead[14]),
        .I1(out[1]),
        .I2(pc_reg[14]_0),
        .I3(memAWrite[14]_i_5_n_0),
        .I4(memAWrite[14]_i_6_n_0),
        .I5(decodedOpcode_reg[3])
    );
    LUT6 memAWrite[14]_i_3
    (
        .O(memAWrite[14]_i_3_n_0),
        .I0(mem_read_IBUF[14]),
        .I1(out[0]),
        .I2(memAWrite_reg[15]_i_5_n_5),
        .I3(out[1]),
        .I4(memBRead[14]),
        .I5(memARead[14])
    );
    LUT6 memAWrite[14]_i_5
    (
        .O(memAWrite[14]_i_5_n_0),
        .I0(memARead[14]),
        .I1(Q[3]),
        .I2(memARead[7]),
        .I3(Q[2]),
        .I4(Q[0]),
        .I5(idim_flag)
    );
    LUT4 memAWrite[14]_i_6
    (
        .O(memAWrite[14]_i_6_n_0),
        .I0(Q[0]),
        .I1(Q[3]),
        .I2(Q[2]),
        .I3(memARead[17])
    );
    LUT6 memAWrite[15]_i_1
    (
        .O(memAWrite_reg[31][15]),
        .I0(memBRead[15]),
        .I1(out[3]),
        .I2(memAWrite[15]_i_2_n_0),
        .I3(out[1]),
        .I4(out[2]),
        .I5(memAWrite[15]_i_3_n_0)
    );
    LUT6 memAWrite[15]_i_2
    (
        .O(memAWrite[15]_i_2_n_0),
        .I0(out[1]),
        .I1(decodedOpcode_reg[2]_0),
        .I2(memARead[15]),
        .I3(decodedOpcode_reg[2]),
        .I4(memARead[16]),
        .I5(memAWrite[15]_i_4_n_0)
    );
    LUT6 memAWrite[15]_i_3
    (
        .O(memAWrite[15]_i_3_n_0),
        .I0(mem_read_IBUF[15]),
        .I1(out[0]),
        .I2(memAWrite_reg[15]_i_5_n_4),
        .I3(out[1]),
        .I4(memBRead[15]),
        .I5(memARead[15])
    );
    LUT5 memAWrite[15]_i_4
    (
        .O(memAWrite[15]_i_4_n_0),
        .I0(memARead[8]),
        .I1(idim_flag),
        .I2(opcode_reg[6]_0[4]),
        .I3(Q[0]),
        .I4(Q[2])
    );
    LUT2 memAWrite[15]_i_6
    (
        .O(memAWrite[15]_i_6_n_0),
        .I0(memARead[15]),
        .I1(memBRead[15])
    );
    LUT2 memAWrite[15]_i_7
    (
        .O(memAWrite[15]_i_7_n_0),
        .I0(memARead[14]),
        .I1(memBRead[14])
    );
    LUT2 memAWrite[15]_i_8
    (
        .O(memAWrite[15]_i_8_n_0),
        .I0(memARead[13]),
        .I1(memBRead[13])
    );
    LUT2 memAWrite[15]_i_9
    (
        .O(memAWrite[15]_i_9_n_0),
        .I0(memARead[12]),
        .I1(memBRead[12])
    );
    LUT6 memAWrite[16]_i_1
    (
        .O(memAWrite_reg[31][16]),
        .I0(memBRead[16]),
        .I1(out[3]),
        .I2(memAWrite[16]_i_2_n_0),
        .I3(out[1]),
        .I4(out[2]),
        .I5(memAWrite[16]_i_3_n_0)
    );
    LUT6 memAWrite[16]_i_2
    (
        .O(memAWrite[16]_i_2_n_0),
        .I0(out[1]),
        .I1(decodedOpcode_reg[2]_0),
        .I2(memARead[16]),
        .I3(decodedOpcode_reg[2]),
        .I4(memARead[15]),
        .I5(memAWrite[16]_i_4_n_0)
    );
    LUT6 memAWrite[16]_i_3
    (
        .O(memAWrite[16]_i_3_n_0),
        .I0(mem_read_IBUF[16]),
        .I1(out[0]),
        .I2(memAWrite_reg[19]_i_5_n_7),
        .I3(out[1]),
        .I4(memBRead[16]),
        .I5(memARead[16])
    );
    LUT5 memAWrite[16]_i_4
    (
        .O(memAWrite[16]_i_4_n_0),
        .I0(memARead[9]),
        .I1(idim_flag),
        .I2(opcode_reg[6]_0[4]),
        .I3(Q[0]),
        .I4(Q[2])
    );
    LUT6 memAWrite[17]_i_1
    (
        .O(memAWrite_reg[31][17]),
        .I0(memBRead[17]),
        .I1(out[3]),
        .I2(memAWrite[17]_i_2_n_0),
        .I3(out[1]),
        .I4(out[2]),
        .I5(memAWrite[17]_i_3_n_0)
    );
    LUT6 memAWrite[17]_i_2
    (
        .O(memAWrite[17]_i_2_n_0),
        .I0(out[1]),
        .I1(decodedOpcode_reg[2]_0),
        .I2(memARead[17]),
        .I3(decodedOpcode_reg[2]),
        .I4(memARead[14]),
        .I5(memAWrite[17]_i_4_n_0)
    );
    LUT6 memAWrite[17]_i_3
    (
        .O(memAWrite[17]_i_3_n_0),
        .I0(mem_read_IBUF[17]),
        .I1(out[0]),
        .I2(memAWrite_reg[19]_i_5_n_6),
        .I3(out[1]),
        .I4(memBRead[17]),
        .I5(memARead[17])
    );
    LUT5 memAWrite[17]_i_4
    (
        .O(memAWrite[17]_i_4_n_0),
        .I0(memARead[10]),
        .I1(idim_flag),
        .I2(opcode_reg[6]_0[4]),
        .I3(Q[0]),
        .I4(Q[2])
    );
    LUT6 memAWrite[18]_i_1
    (
        .O(memAWrite_reg[31][18]),
        .I0(memBRead[18]),
        .I1(out[3]),
        .I2(memAWrite[18]_i_2_n_0),
        .I3(out[1]),
        .I4(out[2]),
        .I5(memAWrite[18]_i_3_n_0)
    );
    LUT6 memAWrite[18]_i_2
    (
        .O(memAWrite[18]_i_2_n_0),
        .I0(out[1]),
        .I1(decodedOpcode_reg[2]_0),
        .I2(memARead[18]),
        .I3(decodedOpcode_reg[2]),
        .I4(memARead[13]),
        .I5(memAWrite[18]_i_4_n_0)
    );
    LUT6 memAWrite[18]_i_3
    (
        .O(memAWrite[18]_i_3_n_0),
        .I0(mem_read_IBUF[18]),
        .I1(out[0]),
        .I2(memAWrite_reg[19]_i_5_n_5),
        .I3(out[1]),
        .I4(memBRead[18]),
        .I5(memARead[18])
    );
    LUT5 memAWrite[18]_i_4
    (
        .O(memAWrite[18]_i_4_n_0),
        .I0(memARead[11]),
        .I1(idim_flag),
        .I2(opcode_reg[6]_0[4]),
        .I3(Q[0]),
        .I4(Q[2])
    );
    LUT6 memAWrite[19]_i_1
    (
        .O(memAWrite_reg[31][19]),
        .I0(memBRead[19]),
        .I1(out[3]),
        .I2(memAWrite[19]_i_2_n_0),
        .I3(out[1]),
        .I4(out[2]),
        .I5(memAWrite[19]_i_3_n_0)
    );
    LUT6 memAWrite[19]_i_2
    (
        .O(memAWrite[19]_i_2_n_0),
        .I0(out[1]),
        .I1(decodedOpcode_reg[2]_0),
        .I2(memARead[19]),
        .I3(decodedOpcode_reg[2]),
        .I4(memARead[12]),
        .I5(memAWrite[19]_i_4_n_0)
    );
    LUT6 memAWrite[19]_i_3
    (
        .O(memAWrite[19]_i_3_n_0),
        .I0(mem_read_IBUF[19]),
        .I1(out[0]),
        .I2(memAWrite_reg[19]_i_5_n_4),
        .I3(out[1]),
        .I4(memBRead[19]),
        .I5(memARead[19])
    );
    LUT5 memAWrite[19]_i_4
    (
        .O(memAWrite[19]_i_4_n_0),
        .I0(memARead[12]),
        .I1(idim_flag),
        .I2(opcode_reg[6]_0[4]),
        .I3(Q[0]),
        .I4(Q[2])
    );
    LUT2 memAWrite[19]_i_6
    (
        .O(memAWrite[19]_i_6_n_0),
        .I0(memARead[19]),
        .I1(memBRead[19])
    );
    LUT2 memAWrite[19]_i_7
    (
        .O(memAWrite[19]_i_7_n_0),
        .I0(memARead[18]),
        .I1(memBRead[18])
    );
    LUT2 memAWrite[19]_i_8
    (
        .O(memAWrite[19]_i_8_n_0),
        .I0(memARead[17]),
        .I1(memBRead[17])
    );
    LUT2 memAWrite[19]_i_9
    (
        .O(memAWrite[19]_i_9_n_0),
        .I0(memARead[16]),
        .I1(memBRead[16])
    );
    LUT6 memAWrite[1]_i_1
    (
        .O(memAWrite_reg[31][1]),
        .I0(memBRead[1]),
        .I1(out[3]),
        .I2(memAWrite[1]_i_2_n_0),
        .I3(out[1]),
        .I4(out[2]),
        .I5(memAWrite[1]_i_3_n_0)
    );
    LUT6 memAWrite[1]_i_2
    (
        .O(memAWrite[1]_i_2_n_0),
        .I0(memARead[1]),
        .I1(out[1]),
        .I2(decodedOpcode_reg[2]),
        .I3(memARead[30]),
        .I4(opcode_reg[1]_0),
        .I5(memAWrite[1]_i_5_n_0)
    );
    LUT6 memAWrite[1]_i_3
    (
        .O(memAWrite[1]_i_3_n_0),
        .I0(mem_read_IBUF[1]),
        .I1(out[0]),
        .I2(memAWrite_reg[3]_i_7_n_6),
        .I3(out[1]),
        .I4(memBRead[1]),
        .I5(memARead[1])
    );
    LUT5 memAWrite[1]_i_5
    (
        .O(memAWrite[1]_i_5_n_0),
        .I0(memARead[1]),
        .I1(Q[0]),
        .I2(pc_reg[14]_1[0]),
        .I3(Q[2]),
        .I4(Q[3])
    );
    LUT6 memAWrite[20]_i_1
    (
        .O(memAWrite_reg[31][20]),
        .I0(memBRead[20]),
        .I1(out[3]),
        .I2(memAWrite[20]_i_2_n_0),
        .I3(out[1]),
        .I4(out[2]),
        .I5(memAWrite[20]_i_3_n_0)
    );
    LUT6 memAWrite[20]_i_2
    (
        .O(memAWrite[20]_i_2_n_0),
        .I0(out[1]),
        .I1(decodedOpcode_reg[2]_0),
        .I2(memARead[20]),
        .I3(decodedOpcode_reg[2]),
        .I4(memARead[11]),
        .I5(memAWrite[20]_i_4_n_0)
    );
    LUT6 memAWrite[20]_i_3
    (
        .O(memAWrite[20]_i_3_n_0),
        .I0(mem_read_IBUF[20]),
        .I1(out[0]),
        .I2(memAWrite_reg[23]_i_5_n_7),
        .I3(out[1]),
        .I4(memBRead[20]),
        .I5(memARead[20])
    );
    LUT5 memAWrite[20]_i_4
    (
        .O(memAWrite[20]_i_4_n_0),
        .I0(memARead[13]),
        .I1(idim_flag),
        .I2(opcode_reg[6]_0[4]),
        .I3(Q[0]),
        .I4(Q[2])
    );
    LUT6 memAWrite[21]_i_1
    (
        .O(memAWrite_reg[31][21]),
        .I0(memBRead[21]),
        .I1(out[3]),
        .I2(memAWrite[21]_i_2_n_0),
        .I3(out[1]),
        .I4(out[2]),
        .I5(memAWrite[21]_i_3_n_0)
    );
    LUT6 memAWrite[21]_i_2
    (
        .O(memAWrite[21]_i_2_n_0),
        .I0(out[1]),
        .I1(decodedOpcode_reg[2]_0),
        .I2(memARead[21]),
        .I3(decodedOpcode_reg[2]),
        .I4(memARead[10]),
        .I5(memAWrite[21]_i_4_n_0)
    );
    LUT6 memAWrite[21]_i_3
    (
        .O(memAWrite[21]_i_3_n_0),
        .I0(mem_read_IBUF[21]),
        .I1(out[0]),
        .I2(memAWrite_reg[23]_i_5_n_6),
        .I3(out[1]),
        .I4(memBRead[21]),
        .I5(memARead[21])
    );
    LUT5 memAWrite[21]_i_4
    (
        .O(memAWrite[21]_i_4_n_0),
        .I0(memARead[14]),
        .I1(idim_flag),
        .I2(opcode_reg[6]_0[4]),
        .I3(Q[0]),
        .I4(Q[2])
    );
    LUT6 memAWrite[22]_i_1
    (
        .O(memAWrite_reg[31][22]),
        .I0(memBRead[22]),
        .I1(out[3]),
        .I2(memAWrite[22]_i_2_n_0),
        .I3(out[1]),
        .I4(out[2]),
        .I5(memAWrite[22]_i_3_n_0)
    );
    LUT6 memAWrite[22]_i_2
    (
        .O(memAWrite[22]_i_2_n_0),
        .I0(out[1]),
        .I1(decodedOpcode_reg[2]_0),
        .I2(memARead[22]),
        .I3(decodedOpcode_reg[2]),
        .I4(memARead[9]),
        .I5(memAWrite[22]_i_4_n_0)
    );
    LUT6 memAWrite[22]_i_3
    (
        .O(memAWrite[22]_i_3_n_0),
        .I0(mem_read_IBUF[22]),
        .I1(out[0]),
        .I2(memAWrite_reg[23]_i_5_n_5),
        .I3(out[1]),
        .I4(memBRead[22]),
        .I5(memARead[22])
    );
    LUT5 memAWrite[22]_i_4
    (
        .O(memAWrite[22]_i_4_n_0),
        .I0(memARead[15]),
        .I1(idim_flag),
        .I2(opcode_reg[6]_0[4]),
        .I3(Q[0]),
        .I4(Q[2])
    );
    LUT6 memAWrite[23]_i_1
    (
        .O(memAWrite_reg[31][23]),
        .I0(memBRead[23]),
        .I1(out[3]),
        .I2(memAWrite[23]_i_2_n_0),
        .I3(out[1]),
        .I4(out[2]),
        .I5(memAWrite[23]_i_3_n_0)
    );
    LUT6 memAWrite[23]_i_2
    (
        .O(memAWrite[23]_i_2_n_0),
        .I0(out[1]),
        .I1(decodedOpcode_reg[2]_0),
        .I2(memARead[23]),
        .I3(decodedOpcode_reg[2]),
        .I4(memARead[8]),
        .I5(memAWrite[23]_i_4_n_0)
    );
    LUT6 memAWrite[23]_i_3
    (
        .O(memAWrite[23]_i_3_n_0),
        .I0(mem_read_IBUF[23]),
        .I1(out[0]),
        .I2(memAWrite_reg[23]_i_5_n_4),
        .I3(out[1]),
        .I4(memBRead[23]),
        .I5(memARead[23])
    );
    LUT5 memAWrite[23]_i_4
    (
        .O(memAWrite[23]_i_4_n_0),
        .I0(memARead[16]),
        .I1(idim_flag),
        .I2(opcode_reg[6]_0[4]),
        .I3(Q[0]),
        .I4(Q[2])
    );
    LUT2 memAWrite[23]_i_6
    (
        .O(memAWrite[23]_i_6_n_0),
        .I0(memARead[23]),
        .I1(memBRead[23])
    );
    LUT2 memAWrite[23]_i_7
    (
        .O(memAWrite[23]_i_7_n_0),
        .I0(memARead[22]),
        .I1(memBRead[22])
    );
    LUT2 memAWrite[23]_i_8
    (
        .O(memAWrite[23]_i_8_n_0),
        .I0(memARead[21]),
        .I1(memBRead[21])
    );
    LUT2 memAWrite[23]_i_9
    (
        .O(memAWrite[23]_i_9_n_0),
        .I0(memARead[20]),
        .I1(memBRead[20])
    );
    LUT6 memAWrite[24]_i_1
    (
        .O(memAWrite_reg[31][24]),
        .I0(memBRead[24]),
        .I1(out[3]),
        .I2(memAWrite[24]_i_2_n_0),
        .I3(out[1]),
        .I4(out[2]),
        .I5(memAWrite[24]_i_3_n_0)
    );
    LUT6 memAWrite[24]_i_2
    (
        .O(memAWrite[24]_i_2_n_0),
        .I0(out[1]),
        .I1(decodedOpcode_reg[2]_0),
        .I2(memARead[24]),
        .I3(decodedOpcode_reg[2]),
        .I4(memARead[7]),
        .I5(memAWrite[24]_i_4_n_0)
    );
    LUT6 memAWrite[24]_i_3
    (
        .O(memAWrite[24]_i_3_n_0),
        .I0(mem_read_IBUF[24]),
        .I1(out[0]),
        .I2(memAWrite_reg[27]_i_5_n_7),
        .I3(out[1]),
        .I4(memBRead[24]),
        .I5(memARead[24])
    );
    LUT5 memAWrite[24]_i_4
    (
        .O(memAWrite[24]_i_4_n_0),
        .I0(memARead[17]),
        .I1(idim_flag),
        .I2(opcode_reg[6]_0[4]),
        .I3(Q[0]),
        .I4(Q[2])
    );
    LUT6 memAWrite[25]_i_1
    (
        .O(memAWrite_reg[31][25]),
        .I0(memBRead[25]),
        .I1(out[3]),
        .I2(memAWrite[25]_i_2_n_0),
        .I3(out[1]),
        .I4(out[2]),
        .I5(memAWrite[25]_i_3_n_0)
    );
    LUT6 memAWrite[25]_i_2
    (
        .O(memAWrite[25]_i_2_n_0),
        .I0(out[1]),
        .I1(decodedOpcode_reg[2]_0),
        .I2(memARead[25]),
        .I3(decodedOpcode_reg[2]),
        .I4(memARead[6]),
        .I5(memAWrite[25]_i_4_n_0)
    );
    LUT6 memAWrite[25]_i_3
    (
        .O(memAWrite[25]_i_3_n_0),
        .I0(mem_read_IBUF[25]),
        .I1(out[0]),
        .I2(memAWrite_reg[27]_i_5_n_6),
        .I3(out[1]),
        .I4(memBRead[25]),
        .I5(memARead[25])
    );
    LUT5 memAWrite[25]_i_4
    (
        .O(memAWrite[25]_i_4_n_0),
        .I0(memARead[18]),
        .I1(idim_flag),
        .I2(opcode_reg[6]_0[4]),
        .I3(Q[0]),
        .I4(Q[2])
    );
    LUT6 memAWrite[26]_i_1
    (
        .O(memAWrite_reg[31][26]),
        .I0(memBRead[26]),
        .I1(out[3]),
        .I2(memAWrite[26]_i_2_n_0),
        .I3(out[1]),
        .I4(out[2]),
        .I5(memAWrite[26]_i_3_n_0)
    );
    LUT6 memAWrite[26]_i_2
    (
        .O(memAWrite[26]_i_2_n_0),
        .I0(out[1]),
        .I1(decodedOpcode_reg[2]_0),
        .I2(memARead[26]),
        .I3(decodedOpcode_reg[2]),
        .I4(memARead[5]),
        .I5(memAWrite[26]_i_4_n_0)
    );
    LUT6 memAWrite[26]_i_3
    (
        .O(memAWrite[26]_i_3_n_0),
        .I0(mem_read_IBUF[26]),
        .I1(out[0]),
        .I2(memAWrite_reg[27]_i_5_n_5),
        .I3(out[1]),
        .I4(memBRead[26]),
        .I5(memARead[26])
    );
    LUT5 memAWrite[26]_i_4
    (
        .O(memAWrite[26]_i_4_n_0),
        .I0(memARead[19]),
        .I1(idim_flag),
        .I2(opcode_reg[6]_0[4]),
        .I3(Q[0]),
        .I4(Q[2])
    );
    LUT6 memAWrite[27]_i_1
    (
        .O(memAWrite_reg[31][27]),
        .I0(memBRead[27]),
        .I1(out[3]),
        .I2(memAWrite[27]_i_2_n_0),
        .I3(out[1]),
        .I4(out[2]),
        .I5(memAWrite[27]_i_3_n_0)
    );
    LUT6 memAWrite[27]_i_2
    (
        .O(memAWrite[27]_i_2_n_0),
        .I0(out[1]),
        .I1(decodedOpcode_reg[2]_0),
        .I2(memARead[27]),
        .I3(decodedOpcode_reg[2]),
        .I4(memARead[4]),
        .I5(memAWrite[27]_i_4_n_0)
    );
    LUT6 memAWrite[27]_i_3
    (
        .O(memAWrite[27]_i_3_n_0),
        .I0(mem_read_IBUF[27]),
        .I1(out[0]),
        .I2(memAWrite_reg[27]_i_5_n_4),
        .I3(out[1]),
        .I4(memBRead[27]),
        .I5(memARead[27])
    );
    LUT5 memAWrite[27]_i_4
    (
        .O(memAWrite[27]_i_4_n_0),
        .I0(memARead[20]),
        .I1(idim_flag),
        .I2(opcode_reg[6]_0[4]),
        .I3(Q[0]),
        .I4(Q[2])
    );
    LUT2 memAWrite[27]_i_6
    (
        .O(memAWrite[27]_i_6_n_0),
        .I0(memARead[27]),
        .I1(memBRead[27])
    );
    LUT2 memAWrite[27]_i_7
    (
        .O(memAWrite[27]_i_7_n_0),
        .I0(memARead[26]),
        .I1(memBRead[26])
    );
    LUT2 memAWrite[27]_i_8
    (
        .O(memAWrite[27]_i_8_n_0),
        .I0(memARead[25]),
        .I1(memBRead[25])
    );
    LUT2 memAWrite[27]_i_9
    (
        .O(memAWrite[27]_i_9_n_0),
        .I0(memARead[24]),
        .I1(memBRead[24])
    );
    LUT6 memAWrite[28]_i_1
    (
        .O(memAWrite_reg[31][28]),
        .I0(memBRead[28]),
        .I1(out[3]),
        .I2(memAWrite[28]_i_2_n_0),
        .I3(out[1]),
        .I4(out[2]),
        .I5(memAWrite[28]_i_3_n_0)
    );
    LUT6 memAWrite[28]_i_2
    (
        .O(memAWrite[28]_i_2_n_0),
        .I0(out[1]),
        .I1(decodedOpcode_reg[2]_0),
        .I2(memARead[28]),
        .I3(decodedOpcode_reg[2]),
        .I4(memARead[3]),
        .I5(memAWrite[28]_i_4_n_0)
    );
    LUT6 memAWrite[28]_i_3
    (
        .O(memAWrite[28]_i_3_n_0),
        .I0(mem_read_IBUF[28]),
        .I1(out[0]),
        .I2(memAWrite_reg[31]_i_6_n_7),
        .I3(out[1]),
        .I4(memBRead[28]),
        .I5(memARead[28])
    );
    LUT5 memAWrite[28]_i_4
    (
        .O(memAWrite[28]_i_4_n_0),
        .I0(memARead[21]),
        .I1(idim_flag),
        .I2(opcode_reg[6]_0[4]),
        .I3(Q[0]),
        .I4(Q[2])
    );
    LUT6 memAWrite[29]_i_1
    (
        .O(memAWrite_reg[31][29]),
        .I0(memBRead[29]),
        .I1(out[3]),
        .I2(memAWrite[29]_i_2_n_0),
        .I3(out[1]),
        .I4(out[2]),
        .I5(memAWrite[29]_i_3_n_0)
    );
    LUT6 memAWrite[29]_i_2
    (
        .O(memAWrite[29]_i_2_n_0),
        .I0(out[1]),
        .I1(decodedOpcode_reg[2]_0),
        .I2(memARead[29]),
        .I3(decodedOpcode_reg[2]),
        .I4(memARead[2]),
        .I5(memAWrite[29]_i_4_n_0)
    );
    LUT6 memAWrite[29]_i_3
    (
        .O(memAWrite[29]_i_3_n_0),
        .I0(mem_read_IBUF[29]),
        .I1(out[0]),
        .I2(memAWrite_reg[31]_i_6_n_6),
        .I3(out[1]),
        .I4(memBRead[29]),
        .I5(memARead[29])
    );
    LUT5 memAWrite[29]_i_4
    (
        .O(memAWrite[29]_i_4_n_0),
        .I0(memARead[22]),
        .I1(idim_flag),
        .I2(opcode_reg[6]_0[4]),
        .I3(Q[0]),
        .I4(Q[2])
    );
    LUT6 memAWrite[2]_i_1
    (
        .O(memAWrite_reg[31][2]),
        .I0(memBRead[2]),
        .I1(out[3]),
        .I2(memAWrite[2]_i_2_n_0),
        .I3(out[1]),
        .I4(out[2]),
        .I5(memAWrite[2]_i_3_n_0)
    );
    LUT5 memAWrite[2]_i_2
    (
        .O(memAWrite[2]_i_2_n_0),
        .I0(memARead[2]),
        .I1(out[1]),
        .I2(pc_reg[2]),
        .I3(decodedOpcode_reg[3]_11),
        .I4(memAWrite[2]_i_6_n_0)
    );
    LUT6 memAWrite[2]_i_3
    (
        .O(memAWrite[2]_i_3_n_0),
        .I0(mem_read_IBUF[2]),
        .I1(out[0]),
        .I2(memAWrite_reg[3]_i_7_n_5),
        .I3(out[1]),
        .I4(memBRead[2]),
        .I5(memARead[2])
    );
    LUT5 memAWrite[2]_i_6
    (
        .O(memAWrite[2]_i_6_n_0),
        .I0(memARead[29]),
        .I1(memARead[2]),
        .I2(Q[2]),
        .I3(Q[3]),
        .I4(Q[0])
    );
    LUT6 memAWrite[30]_i_1
    (
        .O(memAWrite_reg[31][30]),
        .I0(memBRead[30]),
        .I1(out[3]),
        .I2(memAWrite[30]_i_2_n_0),
        .I3(out[1]),
        .I4(out[2]),
        .I5(memAWrite[30]_i_3_n_0)
    );
    LUT6 memAWrite[30]_i_2
    (
        .O(memAWrite[30]_i_2_n_0),
        .I0(out[1]),
        .I1(decodedOpcode_reg[2]_0),
        .I2(memARead[30]),
        .I3(decodedOpcode_reg[2]),
        .I4(memARead[1]),
        .I5(memAWrite[30]_i_4_n_0)
    );
    LUT6 memAWrite[30]_i_3
    (
        .O(memAWrite[30]_i_3_n_0),
        .I0(mem_read_IBUF[30]),
        .I1(out[0]),
        .I2(memAWrite_reg[31]_i_6_n_5),
        .I3(out[1]),
        .I4(memBRead[30]),
        .I5(memARead[30])
    );
    LUT5 memAWrite[30]_i_4
    (
        .O(memAWrite[30]_i_4_n_0),
        .I0(memARead[23]),
        .I1(idim_flag),
        .I2(opcode_reg[6]_0[4]),
        .I3(Q[0]),
        .I4(Q[2])
    );
    LUT6 memAWrite[31]_i_1
    (
        .O(memAWrite_reg[31][31]),
        .I0(memBRead[31]),
        .I1(out[3]),
        .I2(memAWrite[31]_i_2_n_0),
        .I3(out[1]),
        .I4(out[2]),
        .I5(memAWrite[31]_i_3_n_0)
    );
    LUT2 memAWrite[31]_i_10
    (
        .O(memAWrite[31]_i_10_n_0),
        .I0(memARead[28]),
        .I1(memBRead[28])
    );
    LUT6 memAWrite[31]_i_2
    (
        .O(memAWrite[31]_i_2_n_0),
        .I0(out[1]),
        .I1(decodedOpcode_reg[2]_0),
        .I2(memARead[31]),
        .I3(decodedOpcode_reg[2]),
        .I4(memARead[0]),
        .I5(memAWrite[31]_i_5_n_0)
    );
    LUT6 memAWrite[31]_i_3
    (
        .O(memAWrite[31]_i_3_n_0),
        .I0(mem_read_IBUF[31]),
        .I1(out[0]),
        .I2(memAWrite_reg[31]_i_6_n_4),
        .I3(out[1]),
        .I4(memBRead[31]),
        .I5(memARead[31])
    );
    LUT5 memAWrite[31]_i_5
    (
        .O(memAWrite[31]_i_5_n_0),
        .I0(memARead[24]),
        .I1(idim_flag),
        .I2(opcode_reg[6]_0[4]),
        .I3(Q[0]),
        .I4(Q[2])
    );
    LUT2 memAWrite[31]_i_7
    (
        .O(memAWrite[31]_i_7_n_0),
        .I0(memARead[31]),
        .I1(memBRead[31])
    );
    LUT2 memAWrite[31]_i_8
    (
        .O(memAWrite[31]_i_8_n_0),
        .I0(memARead[30]),
        .I1(memBRead[30])
    );
    LUT2 memAWrite[31]_i_9
    (
        .O(memAWrite[31]_i_9_n_0),
        .I0(memARead[29]),
        .I1(memBRead[29])
    );
    LUT6 memAWrite[3]_i_1
    (
        .O(memAWrite_reg[31][3]),
        .I0(memBRead[3]),
        .I1(out[3]),
        .I2(memAWrite[3]_i_2_n_0),
        .I3(out[1]),
        .I4(out[2]),
        .I5(memAWrite[3]_i_3_n_0)
    );
    LUT2 memAWrite[3]_i_10
    (
        .O(memAWrite[3]_i_10_n_0),
        .I0(memARead[1]),
        .I1(memBRead[1])
    );
    LUT2 memAWrite[3]_i_11
    (
        .O(memAWrite[3]_i_11_n_0),
        .I0(memARead[0]),
        .I1(memBRead[0])
    );
    LUT5 memAWrite[3]_i_2
    (
        .O(memAWrite[3]_i_2_n_0),
        .I0(memARead[3]),
        .I1(out[1]),
        .I2(pc_reg[3]),
        .I3(decodedOpcode_reg[3]_10),
        .I4(memAWrite[3]_i_6_n_0)
    );
    LUT6 memAWrite[3]_i_3
    (
        .O(memAWrite[3]_i_3_n_0),
        .I0(mem_read_IBUF[3]),
        .I1(out[0]),
        .I2(memAWrite_reg[3]_i_7_n_4),
        .I3(out[1]),
        .I4(memBRead[3]),
        .I5(memARead[3])
    );
    LUT5 memAWrite[3]_i_6
    (
        .O(memAWrite[3]_i_6_n_0),
        .I0(memARead[28]),
        .I1(memARead[3]),
        .I2(Q[2]),
        .I3(Q[3]),
        .I4(Q[0])
    );
    LUT2 memAWrite[3]_i_8
    (
        .O(memAWrite[3]_i_8_n_0),
        .I0(memARead[3]),
        .I1(memBRead[3])
    );
    LUT2 memAWrite[3]_i_9
    (
        .O(memAWrite[3]_i_9_n_0),
        .I0(memARead[2]),
        .I1(memBRead[2])
    );
    LUT6 memAWrite[4]_i_1
    (
        .O(memAWrite_reg[31][4]),
        .I0(memBRead[4]),
        .I1(out[3]),
        .I2(memAWrite[4]_i_2_n_0),
        .I3(out[1]),
        .I4(out[2]),
        .I5(memAWrite[4]_i_3_n_0)
    );
    LUT5 memAWrite[4]_i_2
    (
        .O(memAWrite[4]_i_2_n_0),
        .I0(memARead[4]),
        .I1(out[1]),
        .I2(pc_reg[4]),
        .I3(decodedOpcode_reg[3]_9),
        .I4(memAWrite[4]_i_6_n_0)
    );
    LUT6 memAWrite[4]_i_3
    (
        .O(memAWrite[4]_i_3_n_0),
        .I0(mem_read_IBUF[4]),
        .I1(out[0]),
        .I2(memAWrite_reg[7]_i_8_n_7),
        .I3(out[1]),
        .I4(memBRead[4]),
        .I5(memARead[4])
    );
    LUT5 memAWrite[4]_i_6
    (
        .O(memAWrite[4]_i_6_n_0),
        .I0(memARead[27]),
        .I1(memARead[4]),
        .I2(Q[2]),
        .I3(Q[3]),
        .I4(Q[0])
    );
    LUT6 memAWrite[5]_i_1
    (
        .O(memAWrite_reg[31][5]),
        .I0(memBRead[5]),
        .I1(out[3]),
        .I2(memAWrite[5]_i_2_n_0),
        .I3(out[1]),
        .I4(out[2]),
        .I5(memAWrite[5]_i_3_n_0)
    );
    LUT5 memAWrite[5]_i_2
    (
        .O(memAWrite[5]_i_2_n_0),
        .I0(memARead[5]),
        .I1(out[1]),
        .I2(pc_reg[5]),
        .I3(decodedOpcode_reg[3]_8),
        .I4(memAWrite[5]_i_6_n_0)
    );
    LUT6 memAWrite[5]_i_3
    (
        .O(memAWrite[5]_i_3_n_0),
        .I0(mem_read_IBUF[5]),
        .I1(out[0]),
        .I2(memAWrite_reg[7]_i_8_n_6),
        .I3(out[1]),
        .I4(memBRead[5]),
        .I5(memARead[5])
    );
    LUT5 memAWrite[5]_i_6
    (
        .O(memAWrite[5]_i_6_n_0),
        .I0(memARead[26]),
        .I1(memARead[5]),
        .I2(Q[2]),
        .I3(Q[3]),
        .I4(Q[0])
    );
    LUT6 memAWrite[6]_i_1
    (
        .O(memAWrite_reg[31][6]),
        .I0(memBRead[6]),
        .I1(out[3]),
        .I2(memAWrite[6]_i_2_n_0),
        .I3(out[1]),
        .I4(out[2]),
        .I5(memAWrite[6]_i_3_n_0)
    );
    LUT5 memAWrite[6]_i_2
    (
        .O(memAWrite[6]_i_2_n_0),
        .I0(memARead[6]),
        .I1(out[1]),
        .I2(pc_reg[6]),
        .I3(decodedOpcode_reg[3]_7),
        .I4(memAWrite[6]_i_6_n_0)
    );
    LUT6 memAWrite[6]_i_3
    (
        .O(memAWrite[6]_i_3_n_0),
        .I0(mem_read_IBUF[6]),
        .I1(out[0]),
        .I2(memAWrite_reg[7]_i_8_n_5),
        .I3(out[1]),
        .I4(memBRead[6]),
        .I5(memARead[6])
    );
    LUT5 memAWrite[6]_i_6
    (
        .O(memAWrite[6]_i_6_n_0),
        .I0(memARead[25]),
        .I1(memARead[6]),
        .I2(Q[2]),
        .I3(Q[3]),
        .I4(Q[0])
    );
    LUT6 memAWrite[7]_i_1
    (
        .O(memAWrite_reg[31][7]),
        .I0(memBRead[7]),
        .I1(out[3]),
        .I2(memAWrite[7]_i_2_n_0),
        .I3(out[1]),
        .I4(out[2]),
        .I5(memAWrite[7]_i_3_n_0)
    );
    LUT2 memAWrite[7]_i_10
    (
        .O(memAWrite[7]_i_10_n_0),
        .I0(memARead[6]),
        .I1(memBRead[6])
    );
    LUT2 memAWrite[7]_i_11
    (
        .O(memAWrite[7]_i_11_n_0),
        .I0(memARead[5]),
        .I1(memBRead[5])
    );
    LUT2 memAWrite[7]_i_12
    (
        .O(memAWrite[7]_i_12_n_0),
        .I0(memARead[4]),
        .I1(memBRead[4])
    );
    LUT6 memAWrite[7]_i_2
    (
        .O(memAWrite[7]_i_2_n_0),
        .I0(memARead[7]),
        .I1(out[1]),
        .I2(pc_reg[7]),
        .I3(memAWrite[7]_i_5_n_0),
        .I4(memAWrite[7]_i_6_n_0),
        .I5(decodedOpcode_reg[3]_6)
    );
    LUT6 memAWrite[7]_i_3
    (
        .O(memAWrite[7]_i_3_n_0),
        .I0(mem_read_IBUF[7]),
        .I1(out[0]),
        .I2(memAWrite_reg[7]_i_8_n_4),
        .I3(out[1]),
        .I4(memBRead[7]),
        .I5(memARead[7])
    );
    LUT6 memAWrite[7]_i_5
    (
        .O(memAWrite[7]_i_5_n_0),
        .I0(memARead[7]),
        .I1(Q[3]),
        .I2(memARead[0]),
        .I3(Q[2]),
        .I4(Q[0]),
        .I5(idim_flag)
    );
    LUT4 memAWrite[7]_i_6
    (
        .O(memAWrite[7]_i_6_n_0),
        .I0(Q[0]),
        .I1(Q[3]),
        .I2(Q[2]),
        .I3(memARead[24])
    );
    LUT2 memAWrite[7]_i_9
    (
        .O(memAWrite[7]_i_9_n_0),
        .I0(memARead[7]),
        .I1(memBRead[7])
    );
    LUT6 memAWrite[8]_i_1
    (
        .O(memAWrite_reg[31][8]),
        .I0(memBRead[8]),
        .I1(out[3]),
        .I2(memAWrite[8]_i_2_n_0),
        .I3(out[1]),
        .I4(out[2]),
        .I5(memAWrite[8]_i_3_n_0)
    );
    LUT6 memAWrite[8]_i_2
    (
        .O(memAWrite[8]_i_2_n_0),
        .I0(memARead[8]),
        .I1(out[1]),
        .I2(pc_reg[8]),
        .I3(memAWrite[8]_i_5_n_0),
        .I4(memAWrite[8]_i_6_n_0),
        .I5(decodedOpcode_reg[3]_5)
    );
    LUT6 memAWrite[8]_i_3
    (
        .O(memAWrite[8]_i_3_n_0),
        .I0(mem_read_IBUF[8]),
        .I1(out[0]),
        .I2(memAWrite_reg[11]_i_8_n_7),
        .I3(out[1]),
        .I4(memBRead[8]),
        .I5(memARead[8])
    );
    LUT6 memAWrite[8]_i_5
    (
        .O(memAWrite[8]_i_5_n_0),
        .I0(memARead[8]),
        .I1(Q[3]),
        .I2(memARead[1]),
        .I3(Q[2]),
        .I4(Q[0]),
        .I5(idim_flag)
    );
    LUT4 memAWrite[8]_i_6
    (
        .O(memAWrite[8]_i_6_n_0),
        .I0(Q[0]),
        .I1(Q[3]),
        .I2(Q[2]),
        .I3(memARead[23])
    );
    LUT6 memAWrite[9]_i_1
    (
        .O(memAWrite_reg[31][9]),
        .I0(memBRead[9]),
        .I1(out[3]),
        .I2(memAWrite[9]_i_2_n_0),
        .I3(out[1]),
        .I4(out[2]),
        .I5(memAWrite[9]_i_3_n_0)
    );
    LUT6 memAWrite[9]_i_2
    (
        .O(memAWrite[9]_i_2_n_0),
        .I0(memARead[9]),
        .I1(out[1]),
        .I2(pc_reg[9]),
        .I3(memAWrite[9]_i_5_n_0),
        .I4(memAWrite[9]_i_6_n_0),
        .I5(decodedOpcode_reg[3]_4)
    );
    LUT6 memAWrite[9]_i_3
    (
        .O(memAWrite[9]_i_3_n_0),
        .I0(mem_read_IBUF[9]),
        .I1(out[0]),
        .I2(memAWrite_reg[11]_i_8_n_6),
        .I3(out[1]),
        .I4(memBRead[9]),
        .I5(memARead[9])
    );
    LUT6 memAWrite[9]_i_5
    (
        .O(memAWrite[9]_i_5_n_0),
        .I0(memARead[9]),
        .I1(Q[3]),
        .I2(memARead[2]),
        .I3(Q[2]),
        .I4(Q[0]),
        .I5(idim_flag)
    );
    LUT4 memAWrite[9]_i_6
    (
        .O(memAWrite[9]_i_6_n_0),
        .I0(Q[0]),
        .I1(Q[3]),
        .I2(Q[2]),
        .I3(memARead[22])
    );
    CARRY4 memAWrite_reg[11]_i_8
    (
        .CI(memAWrite_reg[7]_i_8_n_0),
        .CYINIT(<const0>),
        .CO[3:0]({memAWrite_reg[11]_i_8_n_0, memAWrite_reg[11]_i_8_n_1, memAWrite_reg[11]_i_8_n_2, memAWrite_reg[11]_i_8_n_3}),
        .O[3:0]({memAWrite_reg[11]_i_8_n_4, memAWrite_reg[11]_i_8_n_5, memAWrite_reg[11]_i_8_n_6, memAWrite_reg[11]_i_8_n_7}),
        .DI[3:0]({memARead[11], memARead[10], memARead[9], memARead[8]}),
        .S[3:0]({memAWrite[11]_i_9_n_0, memAWrite[11]_i_10_n_0, memAWrite[11]_i_11_n_0, memAWrite[11]_i_12_n_0})
    );
    CARRY4 memAWrite_reg[15]_i_5
    (
        .CI(memAWrite_reg[11]_i_8_n_0),
        .CYINIT(<const0>),
        .CO[3:0]({memAWrite_reg[15]_i_5_n_0, memAWrite_reg[15]_i_5_n_1, memAWrite_reg[15]_i_5_n_2, memAWrite_reg[15]_i_5_n_3}),
        .O[3:0]({memAWrite_reg[15]_i_5_n_4, memAWrite_reg[15]_i_5_n_5, memAWrite_reg[15]_i_5_n_6, memAWrite_reg[15]_i_5_n_7}),
        .DI[3:0]({memARead[15], memARead[14], memARead[13], memARead[12]}),
        .S[3:0]({memAWrite[15]_i_6_n_0, memAWrite[15]_i_7_n_0, memAWrite[15]_i_8_n_0, memAWrite[15]_i_9_n_0})
    );
    CARRY4 memAWrite_reg[19]_i_5
    (
        .CI(memAWrite_reg[15]_i_5_n_0),
        .CYINIT(<const0>),
        .CO[3:0]({memAWrite_reg[19]_i_5_n_0, memAWrite_reg[19]_i_5_n_1, memAWrite_reg[19]_i_5_n_2, memAWrite_reg[19]_i_5_n_3}),
        .O[3:0]({memAWrite_reg[19]_i_5_n_4, memAWrite_reg[19]_i_5_n_5, memAWrite_reg[19]_i_5_n_6, memAWrite_reg[19]_i_5_n_7}),
        .DI[3:0]({memARead[19], memARead[18], memARead[17], memARead[16]}),
        .S[3:0]({memAWrite[19]_i_6_n_0, memAWrite[19]_i_7_n_0, memAWrite[19]_i_8_n_0, memAWrite[19]_i_9_n_0})
    );
    CARRY4 memAWrite_reg[23]_i_5
    (
        .CI(memAWrite_reg[19]_i_5_n_0),
        .CYINIT(<const0>),
        .CO[3:0]({memAWrite_reg[23]_i_5_n_0, memAWrite_reg[23]_i_5_n_1, memAWrite_reg[23]_i_5_n_2, memAWrite_reg[23]_i_5_n_3}),
        .O[3:0]({memAWrite_reg[23]_i_5_n_4, memAWrite_reg[23]_i_5_n_5, memAWrite_reg[23]_i_5_n_6, memAWrite_reg[23]_i_5_n_7}),
        .DI[3:0]({memARead[23], memARead[22], memARead[21], memARead[20]}),
        .S[3:0]({memAWrite[23]_i_6_n_0, memAWrite[23]_i_7_n_0, memAWrite[23]_i_8_n_0, memAWrite[23]_i_9_n_0})
    );
    CARRY4 memAWrite_reg[27]_i_5
    (
        .CI(memAWrite_reg[23]_i_5_n_0),
        .CYINIT(<const0>),
        .CO[3:0]({memAWrite_reg[27]_i_5_n_0, memAWrite_reg[27]_i_5_n_1, memAWrite_reg[27]_i_5_n_2, memAWrite_reg[27]_i_5_n_3}),
        .O[3:0]({memAWrite_reg[27]_i_5_n_4, memAWrite_reg[27]_i_5_n_5, memAWrite_reg[27]_i_5_n_6, memAWrite_reg[27]_i_5_n_7}),
        .DI[3:0]({memARead[27], memARead[26], memARead[25], memARead[24]}),
        .S[3:0]({memAWrite[27]_i_6_n_0, memAWrite[27]_i_7_n_0, memAWrite[27]_i_8_n_0, memAWrite[27]_i_9_n_0})
    );
    CARRY4 memAWrite_reg[31]_i_6
    (
        .CI(memAWrite_reg[27]_i_5_n_0),
        .CYINIT(<const0>),
        .CO[3:0]({}),
        .O[3:0]({memAWrite_reg[31]_i_6_n_4, memAWrite_reg[31]_i_6_n_5, memAWrite_reg[31]_i_6_n_6, memAWrite_reg[31]_i_6_n_7}),
        .DI[3:0]({<const0>, memARead[30], memARead[29], memARead[28]}),
        .S[3:0]({memAWrite[31]_i_7_n_0, memAWrite[31]_i_8_n_0, memAWrite[31]_i_9_n_0, memAWrite[31]_i_10_n_0})
    );
    CARRY4 memAWrite_reg[3]_i_7
    (
        .CI(<const0>),
        .CYINIT(<const0>),
        .CO[3:0]({memAWrite_reg[3]_i_7_n_0, memAWrite_reg[3]_i_7_n_1, memAWrite_reg[3]_i_7_n_2, memAWrite_reg[3]_i_7_n_3}),
        .O[3:0]({memAWrite_reg[3]_i_7_n_4, memAWrite_reg[3]_i_7_n_5, memAWrite_reg[3]_i_7_n_6, memAWrite_reg[3]_i_7_n_7}),
        .DI[3:0]({memARead[3], memARead[2], memARead[1], memARead[0]}),
        .S[3:0]({memAWrite[3]_i_8_n_0, memAWrite[3]_i_9_n_0, memAWrite[3]_i_10_n_0, memAWrite[3]_i_11_n_0})
    );
    CARRY4 memAWrite_reg[7]_i_8
    (
        .CI(memAWrite_reg[3]_i_7_n_0),
        .CYINIT(<const0>),
        .CO[3:0]({memAWrite_reg[7]_i_8_n_0, memAWrite_reg[7]_i_8_n_1, memAWrite_reg[7]_i_8_n_2, memAWrite_reg[7]_i_8_n_3}),
        .O[3:0]({memAWrite_reg[7]_i_8_n_4, memAWrite_reg[7]_i_8_n_5, memAWrite_reg[7]_i_8_n_6, memAWrite_reg[7]_i_8_n_7}),
        .DI[3:0]({memARead[7], memARead[6], memARead[5], memARead[4]}),
        .S[3:0]({memAWrite[7]_i_9_n_0, memAWrite[7]_i_10_n_0, memAWrite[7]_i_11_n_0, memAWrite[7]_i_12_n_0})
    );
    LUT6 opcode[0]_i_1
    (
        .O(opcode_reg[0]),
        .I0(memBRead[8]),
        .I1(memBRead[0]),
        .I2(pc_reg[1][1]),
        .I3(pc_reg[1][0]),
        .I4(memBRead[24]),
        .I5(memBRead[16])
    );
    LUT6 opcode[1]_i_1
    (
        .O(opcode_reg[1]),
        .I0(memBRead[9]),
        .I1(memBRead[1]),
        .I2(pc_reg[1][1]),
        .I3(pc_reg[1][0]),
        .I4(memBRead[25]),
        .I5(memBRead[17])
    );
    LUT6 opcode[2]_i_1
    (
        .O(opcode_reg[2]),
        .I0(memBRead[10]),
        .I1(memBRead[2]),
        .I2(pc_reg[1][1]),
        .I3(pc_reg[1][0]),
        .I4(memBRead[26]),
        .I5(memBRead[18])
    );
    LUT6 opcode[3]_i_1
    (
        .O(opcode_reg[3]),
        .I0(memBRead[11]),
        .I1(memBRead[3]),
        .I2(pc_reg[1][1]),
        .I3(pc_reg[1][0]),
        .I4(memBRead[27]),
        .I5(memBRead[19])
    );
    LUT6 opcode[4]_i_1
    (
        .O(opcode_reg[4]),
        .I0(memBRead[12]),
        .I1(memBRead[4]),
        .I2(pc_reg[1][1]),
        .I3(pc_reg[1][0]),
        .I4(memBRead[28]),
        .I5(memBRead[20])
    );
    LUT6 opcode[5]_i_1
    (
        .O(opcode_reg[5]),
        .I0(memBRead[13]),
        .I1(memBRead[5]),
        .I2(pc_reg[1][1]),
        .I3(pc_reg[1][0]),
        .I4(memBRead[29]),
        .I5(memBRead[21])
    );
    LUT6 opcode[6]_i_1
    (
        .O(opcode_reg[6]),
        .I0(memBRead[14]),
        .I1(memBRead[6]),
        .I2(pc_reg[1][1]),
        .I3(pc_reg[1][0]),
        .I4(memBRead[30]),
        .I5(memBRead[22])
    );
    LUT5 out_mem_readEnable_i_1
    (
        .O(out_mem_readEnable_reg),
        .I0(decodedOpcode_reg[2]),
        .I1(memARead[15]),
        .I2(Q[1]),
        .I3(Q[4]),
        .I4(FSM_sequential_state_reg[3])
    );
    LUT4 pc[0]_i_1
    (
        .O(pc_reg[14][0]),
        .I0(memARead[0]),
        .I1(decodedOpcode_reg[2]_4),
        .I2(pc_reg[1][0]),
        .I3(decodedOpcode_reg[0]_2)
    );
    LUT4 pc[10]_i_1
    (
        .O(pc_reg[14][10]),
        .I0(memARead[10]),
        .I1(decodedOpcode_reg[2]_4),
        .I2(pc_reg[14]_1[9]),
        .I3(decodedOpcode_reg[0]_2)
    );
    LUT4 pc[11]_i_1
    (
        .O(pc_reg[14][11]),
        .I0(memARead[11]),
        .I1(decodedOpcode_reg[2]_4),
        .I2(pc_reg[14]_1[10]),
        .I3(decodedOpcode_reg[0]_2)
    );
    LUT4 pc[12]_i_1
    (
        .O(pc_reg[14][12]),
        .I0(memARead[12]),
        .I1(decodedOpcode_reg[2]_4),
        .I2(pc_reg[14]_1[11]),
        .I3(decodedOpcode_reg[0]_2)
    );
    LUT4 pc[13]_i_1
    (
        .O(pc_reg[14][13]),
        .I0(memARead[13]),
        .I1(decodedOpcode_reg[2]_4),
        .I2(pc_reg[14]_1[12]),
        .I3(decodedOpcode_reg[0]_2)
    );
    LUT4 pc[14]_i_2
    (
        .O(pc_reg[14][14]),
        .I0(memARead[14]),
        .I1(decodedOpcode_reg[2]_4),
        .I2(pc_reg[14]_1[13]),
        .I3(decodedOpcode_reg[0]_2)
    );
    LUT4 pc[1]_i_1
    (
        .O(pc_reg[14][1]),
        .I0(memARead[1]),
        .I1(decodedOpcode_reg[2]_4),
        .I2(pc_reg[14]_1[0]),
        .I3(decodedOpcode_reg[0]_2)
    );
    LUT4 pc[2]_i_1
    (
        .O(pc_reg[14][2]),
        .I0(memARead[2]),
        .I1(decodedOpcode_reg[2]_4),
        .I2(pc_reg[14]_1[1]),
        .I3(decodedOpcode_reg[0]_2)
    );
    LUT4 pc[3]_i_1
    (
        .O(pc_reg[14][3]),
        .I0(memARead[3]),
        .I1(decodedOpcode_reg[2]_4),
        .I2(pc_reg[14]_1[2]),
        .I3(decodedOpcode_reg[0]_2)
    );
    LUT4 pc[4]_i_1
    (
        .O(pc_reg[14][4]),
        .I0(memARead[4]),
        .I1(decodedOpcode_reg[2]_4),
        .I2(pc_reg[14]_1[3]),
        .I3(decodedOpcode_reg[0]_2)
    );
    LUT6 pc[5]_i_1
    (
        .O(pc_reg[14][5]),
        .I0(opcode_reg[0]_1),
        .I1(decodedOpcode_reg[2]_3),
        .I2(memARead[5]),
        .I3(Q[0]),
        .I4(decodedOpcode_reg[3]_12),
        .I5(pc_reg[14]_1[4])
    );
    LUT6 pc[6]_i_1
    (
        .O(pc_reg[14][6]),
        .I0(decodedOpcode_reg[0]),
        .I1(pc_reg[14]_1[5]),
        .I2(decodedOpcode_reg[0]_0),
        .I3(memARead[6]),
        .I4(opcode_reg[6]_0[0]),
        .I5(decodedOpcode_reg[0]_1)
    );
    LUT6 pc[7]_i_1
    (
        .O(pc_reg[14][7]),
        .I0(decodedOpcode_reg[0]),
        .I1(pc_reg[14]_1[6]),
        .I2(decodedOpcode_reg[0]_0),
        .I3(memARead[7]),
        .I4(opcode_reg[6]_0[1]),
        .I5(decodedOpcode_reg[0]_1)
    );
    LUT6 pc[8]_i_1
    (
        .O(pc_reg[14][8]),
        .I0(decodedOpcode_reg[0]),
        .I1(pc_reg[14]_1[7]),
        .I2(decodedOpcode_reg[0]_0),
        .I3(memARead[8]),
        .I4(opcode_reg[6]_0[2]),
        .I5(decodedOpcode_reg[0]_1)
    );
    LUT6 pc[9]_i_1
    (
        .O(pc_reg[14][9]),
        .I0(decodedOpcode_reg[0]),
        .I1(pc_reg[14]_1[8]),
        .I2(decodedOpcode_reg[0]_0),
        .I3(memARead[9]),
        .I4(opcode_reg[6]_0[3]),
        .I5(decodedOpcode_reg[0]_1)
    );
    RAMB36E1 ram_reg_0
    (
        .CASCADEOUTA(),
        .CASCADEOUTB(),
        .DBITERR(),
        .SBITERR(),
        .CASCADEINA(<const1>),
        .CASCADEINB(<const1>),
        .CLKARDCLK(clk_IBUF_BUFG),
        .CLKBWRCLK(clk_IBUF_BUFG),
        .ENARDEN(<const1>),
        .ENBWREN(<const1>),
        .INJECTDBITERR(),
        .INJECTSBITERR(),
        .REGCEAREGCE(<const0>),
        .REGCEB(<const0>),
        .RSTRAMARSTRAM(<const0>),
        .RSTRAMB(<const0>),
        .RSTREGARSTREG(<const0>),
        .RSTREGB(<const0>),
        .DOADO[31:0]({}),
        .DOBDO[31:0]({}),
        .DOPADOP[3:0](),
        .DOPBDOP[3:0](),
        .ECCPARITY[7:0](),
        .RDADDRECC[8:0](),
        .ADDRARDADDR[15:0]({<const1>, memAAddr_reg[14]_0[12], memAAddr_reg[14]_0[11], memAAddr_reg[14]_0[10], memAAddr_reg[14]_0[9], memAAddr_reg[14]_0[8], memAAddr_reg[14]_0[7], memAAddr_reg[14]_0[6], memAAddr_reg[14]_0[5], memAAddr_reg[14]_0[4], memAAddr_reg[14]_0[3], memAAddr_reg[14]_0[2], memAAddr_reg[14]_0[1], memAAddr_reg[14]_0[0], <const0>, <const0>}),
        .ADDRBWRADDR[15:0]({<const1>, memBAddr_reg[14][12], memBAddr_reg[14][11], memBAddr_reg[14][10], memBAddr_reg[14][9], memBAddr_reg[14][8], memBAddr_reg[14][7], memBAddr_reg[14][6], memBAddr_reg[14][5], memBAddr_reg[14][4], memBAddr_reg[14][3], memBAddr_reg[14][2], memBAddr_reg[14][1], memBAddr_reg[14][0], <const0>, <const0>}),
        .DIADI[31:0]({<const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, memAWrite_reg[31]_0[3], memAWrite_reg[31]_0[2], memAWrite_reg[31]_0[1], memAWrite_reg[31]_0[0]}),
        .DIBDI[31:0]({<const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, memBWrite_reg[31][3], memBWrite_reg[31][2], memBWrite_reg[31][1], memBWrite_reg[31][0]}),
        .DIPADIP[3:0]({<const0>, <const0>, <const0>, <const0>}),
        .DIPBDIP[3:0]({<const0>, <const0>, <const0>, <const0>}),
        .WEA[3:0]({memAWriteEnable, memAWriteEnable, memAWriteEnable, memAWriteEnable}),
        .WEBWE[7:0]({<const0>, <const0>, <const0>, <const0>, memBWriteEnable, memBWriteEnable, memBWriteEnable, memBWriteEnable})
    );
    RAMB36E1 ram_reg_1
    (
        .CASCADEOUTA(),
        .CASCADEOUTB(),
        .DBITERR(),
        .SBITERR(),
        .CASCADEINA(<const1>),
        .CASCADEINB(<const1>),
        .CLKARDCLK(clk_IBUF_BUFG),
        .CLKBWRCLK(clk_IBUF_BUFG),
        .ENARDEN(<const1>),
        .ENBWREN(<const1>),
        .INJECTDBITERR(),
        .INJECTSBITERR(),
        .REGCEAREGCE(<const0>),
        .REGCEB(<const0>),
        .RSTRAMARSTRAM(<const0>),
        .RSTRAMB(<const0>),
        .RSTREGARSTREG(<const0>),
        .RSTREGB(<const0>),
        .DOADO[31:0]({}),
        .DOBDO[31:0]({}),
        .DOPADOP[3:0](),
        .DOPBDOP[3:0](),
        .ECCPARITY[7:0](),
        .RDADDRECC[8:0](),
        .ADDRARDADDR[15:0]({<const1>, memAAddr_reg[14]_0[12], memAAddr_reg[14]_0[11], memAAddr_reg[14]_0[10], memAAddr_reg[14]_0[9], memAAddr_reg[14]_0[8], memAAddr_reg[14]_0[7], memAAddr_reg[14]_0[6], memAAddr_reg[14]_0[5], memAAddr_reg[14]_0[4], memAAddr_reg[14]_0[3], memAAddr_reg[14]_0[2], memAAddr_reg[14]_0[1], memAAddr_reg[14]_0[0], <const0>, <const0>}),
        .ADDRBWRADDR[15:0]({<const1>, memBAddr_reg[14][12], memBAddr_reg[14][11], memBAddr_reg[14][10], memBAddr_reg[14][9], memBAddr_reg[14][8], memBAddr_reg[14][7], memBAddr_reg[14][6], memBAddr_reg[14][5], memBAddr_reg[14][4], memBAddr_reg[14][3], memBAddr_reg[14][2], memBAddr_reg[14][1], memBAddr_reg[14][0], <const0>, <const0>}),
        .DIADI[31:0]({<const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, memAWrite_reg[31]_0[7], memAWrite_reg[31]_0[6], memAWrite_reg[31]_0[5], memAWrite_reg[31]_0[4]}),
        .DIBDI[31:0]({<const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, memBWrite_reg[31][7], memBWrite_reg[31][6], memBWrite_reg[31][5], memBWrite_reg[31][4]}),
        .DIPADIP[3:0]({<const0>, <const0>, <const0>, <const0>}),
        .DIPBDIP[3:0]({<const0>, <const0>, <const0>, <const0>}),
        .WEA[3:0]({memAWriteEnable, memAWriteEnable, memAWriteEnable, memAWriteEnable}),
        .WEBWE[7:0]({<const0>, <const0>, <const0>, <const0>, memBWriteEnable, memBWriteEnable, memBWriteEnable, memBWriteEnable})
    );
    RAMB36E1 ram_reg_2
    (
        .CASCADEOUTA(),
        .CASCADEOUTB(),
        .DBITERR(),
        .SBITERR(),
        .CASCADEINA(<const1>),
        .CASCADEINB(<const1>),
        .CLKARDCLK(clk_IBUF_BUFG),
        .CLKBWRCLK(clk_IBUF_BUFG),
        .ENARDEN(<const1>),
        .ENBWREN(<const1>),
        .INJECTDBITERR(),
        .INJECTSBITERR(),
        .REGCEAREGCE(<const0>),
        .REGCEB(<const0>),
        .RSTRAMARSTRAM(<const0>),
        .RSTRAMB(<const0>),
        .RSTREGARSTREG(<const0>),
        .RSTREGB(<const0>),
        .DOADO[31:0]({}),
        .DOBDO[31:0]({}),
        .DOPADOP[3:0](),
        .DOPBDOP[3:0](),
        .ECCPARITY[7:0](),
        .RDADDRECC[8:0](),
        .ADDRARDADDR[15:0]({<const1>, memAAddr_reg[14]_0[12], memAAddr_reg[14]_0[11], memAAddr_reg[14]_0[10], memAAddr_reg[14]_0[9], memAAddr_reg[14]_0[8], memAAddr_reg[14]_0[7], memAAddr_reg[14]_0[6], memAAddr_reg[14]_0[5], memAAddr_reg[14]_0[4], memAAddr_reg[14]_0[3], memAAddr_reg[14]_0[2], memAAddr_reg[14]_0[1], memAAddr_reg[14]_0[0], <const0>, <const0>}),
        .ADDRBWRADDR[15:0]({<const1>, memBAddr_reg[14][12], memBAddr_reg[14][11], memBAddr_reg[14][10], memBAddr_reg[14][9], memBAddr_reg[14][8], memBAddr_reg[14][7], memBAddr_reg[14][6], memBAddr_reg[14][5], memBAddr_reg[14][4], memBAddr_reg[14][3], memBAddr_reg[14][2], memBAddr_reg[14][1], memBAddr_reg[14][0], <const0>, <const0>}),
        .DIADI[31:0]({<const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, memAWrite_reg[31]_0[11], memAWrite_reg[31]_0[10], memAWrite_reg[31]_0[9], memAWrite_reg[31]_0[8]}),
        .DIBDI[31:0]({<const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, memBWrite_reg[31][11], memBWrite_reg[31][10], memBWrite_reg[31][9], memBWrite_reg[31][8]}),
        .DIPADIP[3:0]({<const0>, <const0>, <const0>, <const0>}),
        .DIPBDIP[3:0]({<const0>, <const0>, <const0>, <const0>}),
        .WEA[3:0]({memAWriteEnable, memAWriteEnable, memAWriteEnable, memAWriteEnable}),
        .WEBWE[7:0]({<const0>, <const0>, <const0>, <const0>, memBWriteEnable, memBWriteEnable, memBWriteEnable, memBWriteEnable})
    );
    RAMB36E1 ram_reg_3
    (
        .CASCADEOUTA(),
        .CASCADEOUTB(),
        .DBITERR(),
        .SBITERR(),
        .CASCADEINA(<const1>),
        .CASCADEINB(<const1>),
        .CLKARDCLK(clk_IBUF_BUFG),
        .CLKBWRCLK(clk_IBUF_BUFG),
        .ENARDEN(<const1>),
        .ENBWREN(<const1>),
        .INJECTDBITERR(),
        .INJECTSBITERR(),
        .REGCEAREGCE(<const0>),
        .REGCEB(<const0>),
        .RSTRAMARSTRAM(<const0>),
        .RSTRAMB(<const0>),
        .RSTREGARSTREG(<const0>),
        .RSTREGB(<const0>),
        .DOADO[31:0]({}),
        .DOBDO[31:0]({}),
        .DOPADOP[3:0](),
        .DOPBDOP[3:0](),
        .ECCPARITY[7:0](),
        .RDADDRECC[8:0](),
        .ADDRARDADDR[15:0]({<const1>, memAAddr_reg[14]_0[12], memAAddr_reg[14]_0[11], memAAddr_reg[14]_0[10], memAAddr_reg[14]_0[9], memAAddr_reg[14]_0[8], memAAddr_reg[14]_0[7], memAAddr_reg[14]_0[6], memAAddr_reg[14]_0[5], memAAddr_reg[14]_0[4], memAAddr_reg[14]_0[3], memAAddr_reg[14]_0[2], memAAddr_reg[14]_0[1], memAAddr_reg[14]_0[0], <const0>, <const0>}),
        .ADDRBWRADDR[15:0]({<const1>, memBAddr_reg[14][12], memBAddr_reg[14][11], memBAddr_reg[14][10], memBAddr_reg[14][9], memBAddr_reg[14][8], memBAddr_reg[14][7], memBAddr_reg[14][6], memBAddr_reg[14][5], memBAddr_reg[14][4], memBAddr_reg[14][3], memBAddr_reg[14][2], memBAddr_reg[14][1], memBAddr_reg[14][0], <const0>, <const0>}),
        .DIADI[31:0]({<const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, memAWrite_reg[31]_0[15], memAWrite_reg[31]_0[14], memAWrite_reg[31]_0[13], memAWrite_reg[31]_0[12]}),
        .DIBDI[31:0]({<const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, memBWrite_reg[31][15], memBWrite_reg[31][14], memBWrite_reg[31][13], memBWrite_reg[31][12]}),
        .DIPADIP[3:0]({<const0>, <const0>, <const0>, <const0>}),
        .DIPBDIP[3:0]({<const0>, <const0>, <const0>, <const0>}),
        .WEA[3:0]({memAWriteEnable, memAWriteEnable, memAWriteEnable, memAWriteEnable}),
        .WEBWE[7:0]({<const0>, <const0>, <const0>, <const0>, memBWriteEnable, memBWriteEnable, memBWriteEnable, memBWriteEnable})
    );
    RAMB36E1 ram_reg_4
    (
        .CASCADEOUTA(),
        .CASCADEOUTB(),
        .DBITERR(),
        .SBITERR(),
        .CASCADEINA(<const1>),
        .CASCADEINB(<const1>),
        .CLKARDCLK(clk_IBUF_BUFG),
        .CLKBWRCLK(clk_IBUF_BUFG),
        .ENARDEN(<const1>),
        .ENBWREN(<const1>),
        .INJECTDBITERR(),
        .INJECTSBITERR(),
        .REGCEAREGCE(<const0>),
        .REGCEB(<const0>),
        .RSTRAMARSTRAM(<const0>),
        .RSTRAMB(<const0>),
        .RSTREGARSTREG(<const0>),
        .RSTREGB(<const0>),
        .DOADO[31:0]({}),
        .DOBDO[31:0]({}),
        .DOPADOP[3:0](),
        .DOPBDOP[3:0](),
        .ECCPARITY[7:0](),
        .RDADDRECC[8:0](),
        .ADDRARDADDR[15:0]({<const1>, memAAddr_reg[14]_0[12], memAAddr_reg[14]_0[11], memAAddr_reg[14]_0[10], memAAddr_reg[14]_0[9], memAAddr_reg[14]_0[8], memAAddr_reg[14]_0[7], memAAddr_reg[14]_0[6], memAAddr_reg[14]_0[5], memAAddr_reg[14]_0[4], memAAddr_reg[14]_0[3], memAAddr_reg[14]_0[2], memAAddr_reg[14]_0[1], memAAddr_reg[14]_0[0], <const0>, <const0>}),
        .ADDRBWRADDR[15:0]({<const1>, memBAddr_reg[14][12], memBAddr_reg[14][11], memBAddr_reg[14][10], memBAddr_reg[14][9], memBAddr_reg[14][8], memBAddr_reg[14][7], memBAddr_reg[14][6], memBAddr_reg[14][5], memBAddr_reg[14][4], memBAddr_reg[14][3], memBAddr_reg[14][2], memBAddr_reg[14][1], memBAddr_reg[14][0], <const0>, <const0>}),
        .DIADI[31:0]({<const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, memAWrite_reg[31]_0[19], memAWrite_reg[31]_0[18], memAWrite_reg[31]_0[17], memAWrite_reg[31]_0[16]}),
        .DIBDI[31:0]({<const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, memBWrite_reg[31][19], memBWrite_reg[31][18], memBWrite_reg[31][17], memBWrite_reg[31][16]}),
        .DIPADIP[3:0]({<const0>, <const0>, <const0>, <const0>}),
        .DIPBDIP[3:0]({<const0>, <const0>, <const0>, <const0>}),
        .WEA[3:0]({memAWriteEnable, memAWriteEnable, memAWriteEnable, memAWriteEnable}),
        .WEBWE[7:0]({<const0>, <const0>, <const0>, <const0>, memBWriteEnable, memBWriteEnable, memBWriteEnable, memBWriteEnable})
    );
    RAMB36E1 ram_reg_5
    (
        .CASCADEOUTA(),
        .CASCADEOUTB(),
        .DBITERR(),
        .SBITERR(),
        .CASCADEINA(<const1>),
        .CASCADEINB(<const1>),
        .CLKARDCLK(clk_IBUF_BUFG),
        .CLKBWRCLK(clk_IBUF_BUFG),
        .ENARDEN(<const1>),
        .ENBWREN(<const1>),
        .INJECTDBITERR(),
        .INJECTSBITERR(),
        .REGCEAREGCE(<const0>),
        .REGCEB(<const0>),
        .RSTRAMARSTRAM(<const0>),
        .RSTRAMB(<const0>),
        .RSTREGARSTREG(<const0>),
        .RSTREGB(<const0>),
        .DOADO[31:0]({}),
        .DOBDO[31:0]({}),
        .DOPADOP[3:0](),
        .DOPBDOP[3:0](),
        .ECCPARITY[7:0](),
        .RDADDRECC[8:0](),
        .ADDRARDADDR[15:0]({<const1>, memAAddr_reg[14]_0[12], memAAddr_reg[14]_0[11], memAAddr_reg[14]_0[10], memAAddr_reg[14]_0[9], memAAddr_reg[14]_0[8], memAAddr_reg[14]_0[7], memAAddr_reg[14]_0[6], memAAddr_reg[14]_0[5], memAAddr_reg[14]_0[4], memAAddr_reg[14]_0[3], memAAddr_reg[14]_0[2], memAAddr_reg[14]_0[1], memAAddr_reg[14]_0[0], <const0>, <const0>}),
        .ADDRBWRADDR[15:0]({<const1>, memBAddr_reg[14][12], memBAddr_reg[14][11], memBAddr_reg[14][10], memBAddr_reg[14][9], memBAddr_reg[14][8], memBAddr_reg[14][7], memBAddr_reg[14][6], memBAddr_reg[14][5], memBAddr_reg[14][4], memBAddr_reg[14][3], memBAddr_reg[14][2], memBAddr_reg[14][1], memBAddr_reg[14][0], <const0>, <const0>}),
        .DIADI[31:0]({<const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, memAWrite_reg[31]_0[23], memAWrite_reg[31]_0[22], memAWrite_reg[31]_0[21], memAWrite_reg[31]_0[20]}),
        .DIBDI[31:0]({<const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, memBWrite_reg[31][23], memBWrite_reg[31][22], memBWrite_reg[31][21], memBWrite_reg[31][20]}),
        .DIPADIP[3:0]({<const0>, <const0>, <const0>, <const0>}),
        .DIPBDIP[3:0]({<const0>, <const0>, <const0>, <const0>}),
        .WEA[3:0]({memAWriteEnable, memAWriteEnable, memAWriteEnable, memAWriteEnable}),
        .WEBWE[7:0]({<const0>, <const0>, <const0>, <const0>, memBWriteEnable, memBWriteEnable, memBWriteEnable, memBWriteEnable})
    );
    RAMB36E1 ram_reg_6
    (
        .CASCADEOUTA(),
        .CASCADEOUTB(),
        .DBITERR(),
        .SBITERR(),
        .CASCADEINA(<const1>),
        .CASCADEINB(<const1>),
        .CLKARDCLK(clk_IBUF_BUFG),
        .CLKBWRCLK(clk_IBUF_BUFG),
        .ENARDEN(<const1>),
        .ENBWREN(<const1>),
        .INJECTDBITERR(),
        .INJECTSBITERR(),
        .REGCEAREGCE(<const0>),
        .REGCEB(<const0>),
        .RSTRAMARSTRAM(<const0>),
        .RSTRAMB(<const0>),
        .RSTREGARSTREG(<const0>),
        .RSTREGB(<const0>),
        .DOADO[31:0]({}),
        .DOBDO[31:0]({}),
        .DOPADOP[3:0](),
        .DOPBDOP[3:0](),
        .ECCPARITY[7:0](),
        .RDADDRECC[8:0](),
        .ADDRARDADDR[15:0]({<const1>, memAAddr_reg[14]_0[12], memAAddr_reg[14]_0[11], memAAddr_reg[14]_0[10], memAAddr_reg[14]_0[9], memAAddr_reg[14]_0[8], memAAddr_reg[14]_0[7], memAAddr_reg[14]_0[6], memAAddr_reg[14]_0[5], memAAddr_reg[14]_0[4], memAAddr_reg[14]_0[3], memAAddr_reg[14]_0[2], memAAddr_reg[14]_0[1], memAAddr_reg[14]_0[0], <const0>, <const0>}),
        .ADDRBWRADDR[15:0]({<const1>, memBAddr_reg[14][12], memBAddr_reg[14][11], memBAddr_reg[14][10], memBAddr_reg[14][9], memBAddr_reg[14][8], memBAddr_reg[14][7], memBAddr_reg[14][6], memBAddr_reg[14][5], memBAddr_reg[14][4], memBAddr_reg[14][3], memBAddr_reg[14][2], memBAddr_reg[14][1], memBAddr_reg[14][0], <const0>, <const0>}),
        .DIADI[31:0]({<const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, memAWrite_reg[31]_0[27], memAWrite_reg[31]_0[26], memAWrite_reg[31]_0[25], memAWrite_reg[31]_0[24]}),
        .DIBDI[31:0]({<const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, memBWrite_reg[31][27], memBWrite_reg[31][26], memBWrite_reg[31][25], memBWrite_reg[31][24]}),
        .DIPADIP[3:0]({<const0>, <const0>, <const0>, <const0>}),
        .DIPBDIP[3:0]({<const0>, <const0>, <const0>, <const0>}),
        .WEA[3:0]({memAWriteEnable, memAWriteEnable, memAWriteEnable, memAWriteEnable}),
        .WEBWE[7:0]({<const0>, <const0>, <const0>, <const0>, memBWriteEnable, memBWriteEnable, memBWriteEnable, memBWriteEnable})
    );
    RAMB36E1 ram_reg_7
    (
        .CASCADEOUTA(),
        .CASCADEOUTB(),
        .DBITERR(),
        .SBITERR(),
        .CASCADEINA(<const1>),
        .CASCADEINB(<const1>),
        .CLKARDCLK(clk_IBUF_BUFG),
        .CLKBWRCLK(clk_IBUF_BUFG),
        .ENARDEN(<const1>),
        .ENBWREN(<const1>),
        .INJECTDBITERR(),
        .INJECTSBITERR(),
        .REGCEAREGCE(<const0>),
        .REGCEB(<const0>),
        .RSTRAMARSTRAM(<const0>),
        .RSTRAMB(<const0>),
        .RSTREGARSTREG(<const0>),
        .RSTREGB(<const0>),
        .DOADO[31:0]({}),
        .DOBDO[31:0]({}),
        .DOPADOP[3:0](),
        .DOPBDOP[3:0](),
        .ECCPARITY[7:0](),
        .RDADDRECC[8:0](),
        .ADDRARDADDR[15:0]({<const1>, memAAddr_reg[14]_0[12], memAAddr_reg[14]_0[11], memAAddr_reg[14]_0[10], memAAddr_reg[14]_0[9], memAAddr_reg[14]_0[8], memAAddr_reg[14]_0[7], memAAddr_reg[14]_0[6], memAAddr_reg[14]_0[5], memAAddr_reg[14]_0[4], memAAddr_reg[14]_0[3], memAAddr_reg[14]_0[2], memAAddr_reg[14]_0[1], memAAddr_reg[14]_0[0], <const0>, <const0>}),
        .ADDRBWRADDR[15:0]({<const1>, memBAddr_reg[14][12], memBAddr_reg[14][11], memBAddr_reg[14][10], memBAddr_reg[14][9], memBAddr_reg[14][8], memBAddr_reg[14][7], memBAddr_reg[14][6], memBAddr_reg[14][5], memBAddr_reg[14][4], memBAddr_reg[14][3], memBAddr_reg[14][2], memBAddr_reg[14][1], memBAddr_reg[14][0], <const0>, <const0>}),
        .DIADI[31:0]({<const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, memAWrite_reg[31]_0[31], memAWrite_reg[31]_0[30], memAWrite_reg[31]_0[29], memAWrite_reg[31]_0[28]}),
        .DIBDI[31:0]({<const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, <const0>, memBWrite_reg[31][31], memBWrite_reg[31][30], memBWrite_reg[31][29], memBWrite_reg[31][28]}),
        .DIPADIP[3:0]({<const0>, <const0>, <const0>, <const0>}),
        .DIPBDIP[3:0]({<const0>, <const0>, <const0>, <const0>}),
        .WEA[3:0]({memAWriteEnable, memAWriteEnable, memAWriteEnable, memAWriteEnable}),
        .WEBWE[7:0]({<const0>, <const0>, <const0>, <const0>, memBWriteEnable, memBWriteEnable, memBWriteEnable, memBWriteEnable})
    );
    LUT6 sp[10]_i_1
    (
        .O(sp_reg[14][8]),
        .I0(out[0]),
        .I1(sp[10]_i_2_n_0),
        .I2(decodedOpcode_reg[2]_1),
        .I3(data2[7]),
        .I4(decodedOpcode_reg[2]_2),
        .I5(sp_reg[10][3])
    );
    LUT4 sp[10]_i_2
    (
        .O(sp[10]_i_2_n_0),
        .I0(memARead[10]),
        .I1(decodedOpcode_reg[0]_4),
        .I2(sp_reg[14]_0[8]),
        .I3(decodedOpcode_reg[4]_0)
    );
    LUT6 sp[11]_i_1
    (
        .O(sp_reg[14][9]),
        .I0(out[0]),
        .I1(sp[11]_i_2_n_0),
        .I2(decodedOpcode_reg[2]_1),
        .I3(data2[8]),
        .I4(decodedOpcode_reg[2]_2),
        .I5(O[0])
    );
    LUT4 sp[11]_i_2
    (
        .O(sp[11]_i_2_n_0),
        .I0(memARead[11]),
        .I1(decodedOpcode_reg[0]_4),
        .I2(sp_reg[14]_0[9]),
        .I3(decodedOpcode_reg[4]_0)
    );
    LUT6 sp[12]_i_1
    (
        .O(sp_reg[14][10]),
        .I0(out[0]),
        .I1(sp[12]_i_2_n_0),
        .I2(decodedOpcode_reg[2]_1),
        .I3(data2[9]),
        .I4(decodedOpcode_reg[2]_2),
        .I5(O[1])
    );
    LUT4 sp[12]_i_2
    (
        .O(sp[12]_i_2_n_0),
        .I0(memARead[12]),
        .I1(decodedOpcode_reg[0]_4),
        .I2(sp_reg[14]_0[10]),
        .I3(decodedOpcode_reg[4]_0)
    );
    LUT6 sp[13]_i_1
    (
        .O(sp_reg[14][11]),
        .I0(out[0]),
        .I1(sp[13]_i_2_n_0),
        .I2(decodedOpcode_reg[2]_1),
        .I3(data2[10]),
        .I4(decodedOpcode_reg[2]_2),
        .I5(O[2])
    );
    LUT4 sp[13]_i_2
    (
        .O(sp[13]_i_2_n_0),
        .I0(memARead[13]),
        .I1(decodedOpcode_reg[0]_4),
        .I2(sp_reg[14]_0[11]),
        .I3(decodedOpcode_reg[4]_0)
    );
    LUT6 sp[14]_i_2
    (
        .O(sp_reg[14][12]),
        .I0(out[0]),
        .I1(sp[14]_i_3_n_0),
        .I2(decodedOpcode_reg[2]_1),
        .I3(data2[11]),
        .I4(decodedOpcode_reg[2]_2),
        .I5(O[3])
    );
    LUT4 sp[14]_i_3
    (
        .O(sp[14]_i_3_n_0),
        .I0(memARead[14]),
        .I1(decodedOpcode_reg[0]_4),
        .I2(sp_reg[14]_0[12]),
        .I3(decodedOpcode_reg[4]_0)
    );
    LUT6 sp[2]_i_1
    (
        .O(sp_reg[14][0]),
        .I0(out[0]),
        .I1(decodedOpcode_reg[4]_0),
        .I2(sp[2]_i_3_n_0),
        .I3(decodedOpcode_reg[2]_1),
        .I4(sp_reg[14]_0[0]),
        .I5(decodedOpcode_reg[2]_2)
    );
    LUT5 sp[2]_i_3
    (
        .O(sp[2]_i_3_n_0),
        .I0(Q[4]),
        .I1(Q[3]),
        .I2(Q[1]),
        .I3(Q[0]),
        .I4(memARead[2])
    );
    LUT6 sp[3]_i_1
    (
        .O(sp_reg[14][1]),
        .I0(out[0]),
        .I1(sp[3]_i_2_n_0),
        .I2(decodedOpcode_reg[2]_1),
        .I3(data2[0]),
        .I4(decodedOpcode_reg[2]_2),
        .I5(sp_reg[2][0])
    );
    LUT4 sp[3]_i_2
    (
        .O(sp[3]_i_2_n_0),
        .I0(memARead[3]),
        .I1(decodedOpcode_reg[0]_4),
        .I2(sp_reg[14]_0[1]),
        .I3(decodedOpcode_reg[4]_0)
    );
    LUT6 sp[4]_i_1
    (
        .O(sp_reg[14][2]),
        .I0(out[0]),
        .I1(sp[4]_i_2_n_0),
        .I2(decodedOpcode_reg[2]_1),
        .I3(data2[1]),
        .I4(decodedOpcode_reg[2]_2),
        .I5(sp_reg[2][1])
    );
    LUT4 sp[4]_i_2
    (
        .O(sp[4]_i_2_n_0),
        .I0(memARead[4]),
        .I1(decodedOpcode_reg[0]_4),
        .I2(sp_reg[14]_0[2]),
        .I3(decodedOpcode_reg[4]_0)
    );
    LUT6 sp[5]_i_1
    (
        .O(sp_reg[14][3]),
        .I0(out[0]),
        .I1(sp[5]_i_2_n_0),
        .I2(decodedOpcode_reg[2]_1),
        .I3(data2[2]),
        .I4(decodedOpcode_reg[2]_2),
        .I5(sp_reg[2][2])
    );
    LUT4 sp[5]_i_2
    (
        .O(sp[5]_i_2_n_0),
        .I0(memARead[5]),
        .I1(decodedOpcode_reg[0]_4),
        .I2(sp_reg[14]_0[3]),
        .I3(decodedOpcode_reg[4]_0)
    );
    LUT6 sp[6]_i_1
    (
        .O(sp_reg[14][4]),
        .I0(out[0]),
        .I1(sp[6]_i_2_n_0),
        .I2(decodedOpcode_reg[2]_1),
        .I3(data2[3]),
        .I4(decodedOpcode_reg[2]_2),
        .I5(sp_reg[2][3])
    );
    LUT4 sp[6]_i_2
    (
        .O(sp[6]_i_2_n_0),
        .I0(memARead[6]),
        .I1(decodedOpcode_reg[0]_4),
        .I2(sp_reg[14]_0[4]),
        .I3(decodedOpcode_reg[4]_0)
    );
    LUT6 sp[7]_i_1
    (
        .O(sp_reg[14][5]),
        .I0(out[0]),
        .I1(sp[7]_i_2_n_0),
        .I2(decodedOpcode_reg[2]_1),
        .I3(data2[4]),
        .I4(decodedOpcode_reg[2]_2),
        .I5(sp_reg[10][0])
    );
    LUT4 sp[7]_i_2
    (
        .O(sp[7]_i_2_n_0),
        .I0(memARead[7]),
        .I1(decodedOpcode_reg[0]_4),
        .I2(sp_reg[14]_0[5]),
        .I3(decodedOpcode_reg[4]_0)
    );
    LUT6 sp[8]_i_1
    (
        .O(sp_reg[14][6]),
        .I0(out[0]),
        .I1(sp[8]_i_2_n_0),
        .I2(decodedOpcode_reg[2]_1),
        .I3(data2[5]),
        .I4(decodedOpcode_reg[2]_2),
        .I5(sp_reg[10][1])
    );
    LUT4 sp[8]_i_2
    (
        .O(sp[8]_i_2_n_0),
        .I0(memARead[8]),
        .I1(decodedOpcode_reg[0]_4),
        .I2(sp_reg[14]_0[6]),
        .I3(decodedOpcode_reg[4]_0)
    );
    LUT6 sp[9]_i_1
    (
        .O(sp_reg[14][7]),
        .I0(out[0]),
        .I1(sp[9]_i_2_n_0),
        .I2(decodedOpcode_reg[2]_1),
        .I3(data2[6]),
        .I4(decodedOpcode_reg[2]_2),
        .I5(sp_reg[10][2])
    );
    LUT4 sp[9]_i_2
    (
        .O(sp[9]_i_2_n_0),
        .I0(memARead[9]),
        .I1(decodedOpcode_reg[0]_4),
        .I2(sp_reg[14]_0[7]),
        .I3(decodedOpcode_reg[4]_0)
    );
endmodule

module FDPE
(
    Q,
    C,
    CE,
    D,
    PRE
);

    output Q;
    input C;
    input CE;
    input D;
    input PRE;


endmodule

module RAMB36E1
(
    CASCADEOUTA,
    CASCADEOUTB,
    DBITERR,
    SBITERR,
    CASCADEINA,
    CASCADEINB,
    CLKARDCLK,
    CLKBWRCLK,
    ENARDEN,
    ENBWREN,
    INJECTDBITERR,
    INJECTSBITERR,
    REGCEAREGCE,
    REGCEB,
    RSTRAMARSTRAM,
    RSTRAMB,
    RSTREGARSTREG,
    RSTREGB,
    DOADO[31:0],
    DOBDO[31:0],
    DOPADOP[3:0],
    DOPBDOP[3:0],
    ECCPARITY[7:0],
    RDADDRECC[8:0],
    ADDRARDADDR[15:0],
    ADDRBWRADDR[15:0],
    DIADI[31:0],
    DIBDI[31:0],
    DIPADIP[3:0],
    DIPBDIP[3:0],
    WEA[3:0],
    WEBWE[7:0]
);

    output CASCADEOUTA;
    output CASCADEOUTB;
    output DBITERR;
    output SBITERR;
    input CASCADEINA;
    input CASCADEINB;
    input CLKARDCLK;
    input CLKBWRCLK;
    input ENARDEN;
    input ENBWREN;
    input INJECTDBITERR;
    input INJECTSBITERR;
    input REGCEAREGCE;
    input REGCEB;
    input RSTRAMARSTRAM;
    input RSTRAMB;
    input RSTREGARSTREG;
    input RSTREGB;
    output [31:0]DOADO[31:0];
    output [31:0]DOBDO[31:0];
    output [3:0]DOPADOP[3:0];
    output [3:0]DOPBDOP[3:0];
    output [7:0]ECCPARITY[7:0];
    output [8:0]RDADDRECC[8:0];
    input [15:0]ADDRARDADDR[15:0];
    input [15:0]ADDRBWRADDR[15:0];
    input [31:0]DIADI[31:0];
    input [31:0]DIBDI[31:0];
    input [3:0]DIPADIP[3:0];
    input [3:0]DIPBDIP[3:0];
    input [3:0]WEA[3:0];
    input [7:0]WEBWE[7:0];


endmodule

module INV
(
    I,
    O
);

    input I;
    output O;


endmodule

