//Generated from netlist by SpyDrNet
//netlist name: random
`celldefine
module $_DLATCHSR_PPP_
(
    D,
    R,
    S,
    E,
    Q
);

    input D;
    input R;
    input S;
    input E;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DLATCHSR_PPN_
(
    D,
    R,
    S,
    E,
    Q
);

    input D;
    input R;
    input S;
    input E;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DLATCHSR_PNP_
(
    D,
    R,
    S,
    E,
    Q
);

    input D;
    input R;
    input S;
    input E;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DLATCHSR_PNN_
(
    D,
    R,
    S,
    E,
    Q
);

    input D;
    input R;
    input S;
    input E;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DLATCHSR_NPP_
(
    D,
    R,
    S,
    E,
    Q
);

    input D;
    input R;
    input S;
    input E;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DLATCHSR_NPN_
(
    D,
    R,
    S,
    E,
    Q
);

    input D;
    input R;
    input S;
    input E;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DLATCHSR_NNP_
(
    D,
    R,
    S,
    E,
    Q
);

    input D;
    input R;
    input S;
    input E;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DLATCHSR_NNN_
(
    D,
    R,
    S,
    E,
    Q
);

    input D;
    input R;
    input S;
    input E;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DLATCH_PP1_
(
    D,
    R,
    E,
    Q
);

    input D;
    input R;
    input E;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DLATCH_PP0_
(
    D,
    R,
    E,
    Q
);

    input D;
    input R;
    input E;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DLATCH_PN1_
(
    D,
    R,
    E,
    Q
);

    input D;
    input R;
    input E;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DLATCH_PN0_
(
    D,
    R,
    E,
    Q
);

    input D;
    input R;
    input E;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DLATCH_NP1_
(
    D,
    R,
    E,
    Q
);

    input D;
    input R;
    input E;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DLATCH_NP0_
(
    D,
    R,
    E,
    Q
);

    input D;
    input R;
    input E;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DLATCH_NN1_
(
    D,
    R,
    E,
    Q
);

    input D;
    input R;
    input E;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DLATCH_NN0_
(
    D,
    R,
    E,
    Q
);

    input D;
    input R;
    input E;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DLATCH_P_
(
    D,
    E,
    Q
);

    input D;
    input E;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DLATCH_N_
(
    D,
    E,
    Q
);

    input D;
    input E;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_SDFFCE_PP1P_
(
    E,
    D,
    R,
    C,
    Q
);

    input E;
    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_SDFFCE_PP1N_
(
    E,
    D,
    R,
    C,
    Q
);

    input E;
    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_SDFFCE_PP0P_
(
    E,
    D,
    R,
    C,
    Q
);

    input E;
    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_SDFFCE_PP0N_
(
    E,
    D,
    R,
    C,
    Q
);

    input E;
    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_SDFFCE_PN1P_
(
    E,
    D,
    R,
    C,
    Q
);

    input E;
    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_SDFFCE_PN1N_
(
    E,
    D,
    R,
    C,
    Q
);

    input E;
    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_SDFFCE_PN0P_
(
    E,
    D,
    R,
    C,
    Q
);

    input E;
    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_SDFFCE_PN0N_
(
    E,
    D,
    R,
    C,
    Q
);

    input E;
    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_SDFFCE_NP1P_
(
    E,
    D,
    R,
    C,
    Q
);

    input E;
    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_SDFFCE_NP1N_
(
    E,
    D,
    R,
    C,
    Q
);

    input E;
    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_SDFFCE_NP0P_
(
    E,
    D,
    R,
    C,
    Q
);

    input E;
    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_SDFFCE_NP0N_
(
    E,
    D,
    R,
    C,
    Q
);

    input E;
    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_SDFFCE_NN1P_
(
    E,
    D,
    R,
    C,
    Q
);

    input E;
    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_SDFFCE_NN1N_
(
    E,
    D,
    R,
    C,
    Q
);

    input E;
    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_SDFFCE_NN0P_
(
    E,
    D,
    R,
    C,
    Q
);

    input E;
    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_SDFFCE_NN0N_
(
    E,
    D,
    R,
    C,
    Q
);

    input E;
    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_SDFFE_PP1P_
(
    E,
    D,
    R,
    C,
    Q
);

    input E;
    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_SDFFE_PP1N_
(
    E,
    D,
    R,
    C,
    Q
);

    input E;
    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_SDFFE_PP0P_
(
    E,
    D,
    R,
    C,
    Q
);

    input E;
    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_SDFFE_PP0N_
(
    E,
    D,
    R,
    C,
    Q
);

    input E;
    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_SDFFE_PN1P_
(
    E,
    D,
    R,
    C,
    Q
);

    input E;
    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_SDFFE_PN1N_
(
    E,
    D,
    R,
    C,
    Q
);

    input E;
    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_SDFFE_PN0P_
(
    E,
    D,
    R,
    C,
    Q
);

    input E;
    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_SDFFE_PN0N_
(
    E,
    D,
    R,
    C,
    Q
);

    input E;
    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_SDFFE_NP1P_
(
    E,
    D,
    R,
    C,
    Q
);

    input E;
    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_SDFFE_NP1N_
(
    E,
    D,
    R,
    C,
    Q
);

    input E;
    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_SDFFE_NP0P_
(
    E,
    D,
    R,
    C,
    Q
);

    input E;
    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_SDFFE_NP0N_
(
    E,
    D,
    R,
    C,
    Q
);

    input E;
    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_SDFFE_NN1P_
(
    E,
    D,
    R,
    C,
    Q
);

    input E;
    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_SDFFE_NN1N_
(
    E,
    D,
    R,
    C,
    Q
);

    input E;
    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_SDFFE_NN0P_
(
    E,
    D,
    R,
    C,
    Q
);

    input E;
    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_SDFFE_NN0N_
(
    E,
    D,
    R,
    C,
    Q
);

    input E;
    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_SDFF_PP1_
(
    D,
    R,
    C,
    Q
);

    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_SDFF_PP0_
(
    D,
    R,
    C,
    Q
);

    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_SDFF_PN1_
(
    D,
    R,
    C,
    Q
);

    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_SDFF_PN0_
(
    D,
    R,
    C,
    Q
);

    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_SDFF_NP1_
(
    D,
    R,
    C,
    Q
);

    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_SDFF_NP0_
(
    D,
    R,
    C,
    Q
);

    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_SDFF_NN1_
(
    D,
    R,
    C,
    Q
);

    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_SDFF_NN0_
(
    D,
    R,
    C,
    Q
);

    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFFSRE_PPPP_
(
    E,
    D,
    R,
    S,
    C,
    Q
);

    input E;
    input D;
    input R;
    input S;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFFSRE_PPPN_
(
    E,
    D,
    R,
    S,
    C,
    Q
);

    input E;
    input D;
    input R;
    input S;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFFSRE_PPNP_
(
    E,
    D,
    R,
    S,
    C,
    Q
);

    input E;
    input D;
    input R;
    input S;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFFSRE_PPNN_
(
    E,
    D,
    R,
    S,
    C,
    Q
);

    input E;
    input D;
    input R;
    input S;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFFSRE_PNPP_
(
    E,
    D,
    R,
    S,
    C,
    Q
);

    input E;
    input D;
    input R;
    input S;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFFSRE_PNPN_
(
    E,
    D,
    R,
    S,
    C,
    Q
);

    input E;
    input D;
    input R;
    input S;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFFSRE_PNNP_
(
    E,
    D,
    R,
    S,
    C,
    Q
);

    input E;
    input D;
    input R;
    input S;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFFSRE_PNNN_
(
    E,
    D,
    R,
    S,
    C,
    Q
);

    input E;
    input D;
    input R;
    input S;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFFSRE_NPPP_
(
    E,
    D,
    R,
    S,
    C,
    Q
);

    input E;
    input D;
    input R;
    input S;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFFSRE_NPPN_
(
    E,
    D,
    R,
    S,
    C,
    Q
);

    input E;
    input D;
    input R;
    input S;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFFSRE_NPNP_
(
    E,
    D,
    R,
    S,
    C,
    Q
);

    input E;
    input D;
    input R;
    input S;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFFSRE_NPNN_
(
    E,
    D,
    R,
    S,
    C,
    Q
);

    input E;
    input D;
    input R;
    input S;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFFSRE_NNPP_
(
    E,
    D,
    R,
    S,
    C,
    Q
);

    input E;
    input D;
    input R;
    input S;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFFSRE_NNPN_
(
    E,
    D,
    R,
    S,
    C,
    Q
);

    input E;
    input D;
    input R;
    input S;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFFSRE_NNNP_
(
    E,
    D,
    R,
    S,
    C,
    Q
);

    input E;
    input D;
    input R;
    input S;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFFSRE_NNNN_
(
    E,
    D,
    R,
    S,
    C,
    Q
);

    input E;
    input D;
    input R;
    input S;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFFSR_PPP_
(
    D,
    R,
    S,
    C,
    Q
);

    input D;
    input R;
    input S;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFFSR_PPN_
(
    D,
    R,
    S,
    C,
    Q
);

    input D;
    input R;
    input S;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFFSR_PNP_
(
    D,
    R,
    S,
    C,
    Q
);

    input D;
    input R;
    input S;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFFSR_PNN_
(
    D,
    R,
    S,
    C,
    Q
);

    input D;
    input R;
    input S;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFFSR_NPP_
(
    D,
    R,
    S,
    C,
    Q
);

    input D;
    input R;
    input S;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFFSR_NPN_
(
    D,
    R,
    S,
    C,
    Q
);

    input D;
    input R;
    input S;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFFSR_NNP_
(
    D,
    R,
    S,
    C,
    Q
);

    input D;
    input R;
    input S;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFFSR_NNN_
(
    D,
    R,
    S,
    C,
    Q
);

    input D;
    input R;
    input S;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_ALDFFE_PPP_
(
    E,
    D,
    AD,
    L,
    C,
    Q
);

    input E;
    input D;
    input AD;
    input L;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_ALDFFE_PPN_
(
    E,
    D,
    AD,
    L,
    C,
    Q
);

    input E;
    input D;
    input AD;
    input L;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_ALDFFE_PNP_
(
    E,
    D,
    AD,
    L,
    C,
    Q
);

    input E;
    input D;
    input AD;
    input L;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_ALDFFE_PNN_
(
    E,
    D,
    AD,
    L,
    C,
    Q
);

    input E;
    input D;
    input AD;
    input L;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_ALDFFE_NPP_
(
    E,
    D,
    AD,
    L,
    C,
    Q
);

    input E;
    input D;
    input AD;
    input L;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_ALDFFE_NPN_
(
    E,
    D,
    AD,
    L,
    C,
    Q
);

    input E;
    input D;
    input AD;
    input L;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_ALDFFE_NNP_
(
    E,
    D,
    AD,
    L,
    C,
    Q
);

    input E;
    input D;
    input AD;
    input L;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_ALDFFE_NNN_
(
    E,
    D,
    AD,
    L,
    C,
    Q
);

    input E;
    input D;
    input AD;
    input L;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_ALDFF_PP_
(
    D,
    AD,
    L,
    C,
    Q
);

    input D;
    input AD;
    input L;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_ALDFF_PN_
(
    D,
    AD,
    L,
    C,
    Q
);

    input D;
    input AD;
    input L;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_ALDFF_NP_
(
    D,
    AD,
    L,
    C,
    Q
);

    input D;
    input AD;
    input L;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_ALDFF_NN_
(
    D,
    AD,
    L,
    C,
    Q
);

    input D;
    input AD;
    input L;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFFE_PP1P_
(
    E,
    D,
    R,
    C,
    Q
);

    input E;
    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFFE_PP1N_
(
    E,
    D,
    R,
    C,
    Q
);

    input E;
    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFFE_PP0P_
(
    E,
    D,
    R,
    C,
    Q
);

    input E;
    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFFE_PP0N_
(
    E,
    D,
    R,
    C,
    Q
);

    input E;
    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFFE_PN1P_
(
    E,
    D,
    R,
    C,
    Q
);

    input E;
    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFFE_PN1N_
(
    E,
    D,
    R,
    C,
    Q
);

    input E;
    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFFE_PN0P_
(
    E,
    D,
    R,
    C,
    Q
);

    input E;
    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFFE_PN0N_
(
    E,
    D,
    R,
    C,
    Q
);

    input E;
    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFFE_NP1P_
(
    E,
    D,
    R,
    C,
    Q
);

    input E;
    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFFE_NP1N_
(
    E,
    D,
    R,
    C,
    Q
);

    input E;
    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFFE_NP0P_
(
    E,
    D,
    R,
    C,
    Q
);

    input E;
    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFFE_NP0N_
(
    E,
    D,
    R,
    C,
    Q
);

    input E;
    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFFE_NN1P_
(
    E,
    D,
    R,
    C,
    Q
);

    input E;
    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFFE_NN1N_
(
    E,
    D,
    R,
    C,
    Q
);

    input E;
    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFFE_NN0P_
(
    E,
    D,
    R,
    C,
    Q
);

    input E;
    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFFE_NN0N_
(
    E,
    D,
    R,
    C,
    Q
);

    input E;
    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFF_PP1_
(
    D,
    R,
    C,
    Q
);

    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFF_PP0_
(
    D,
    R,
    C,
    Q
);

    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFF_PN1_
(
    D,
    R,
    C,
    Q
);

    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFF_PN0_
(
    D,
    R,
    C,
    Q
);

    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFF_NP1_
(
    D,
    R,
    C,
    Q
);

    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFF_NP0_
(
    D,
    R,
    C,
    Q
);

    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFF_NN1_
(
    D,
    R,
    C,
    Q
);

    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFF_NN0_
(
    D,
    R,
    C,
    Q
);

    input D;
    input R;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFFE_PP_
(
    E,
    D,
    C,
    Q
);

    input E;
    input D;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFFE_PN_
(
    E,
    D,
    C,
    Q
);

    input E;
    input D;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFFE_NP_
(
    E,
    D,
    C,
    Q
);

    input E;
    input D;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFFE_NN_
(
    E,
    D,
    C,
    Q
);

    input E;
    input D;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFF_P_
(
    D,
    C,
    Q
);

    input D;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_DFF_N_
(
    D,
    C,
    Q
);

    input D;
    input C;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_FF_
(
    D,
    Q
);

    input D;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_SR_PP_
(
    R,
    S,
    Q
);

    input R;
    input S;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_SR_PN_
(
    R,
    S,
    Q
);

    input R;
    input S;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_SR_NP_
(
    R,
    S,
    Q
);

    input R;
    input S;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_SR_NN_
(
    R,
    S,
    Q
);

    input R;
    input S;
    output Q;

endmodule
`endcelldefine

`celldefine
module $_TBUF_
(
    E,
    A,
    Y
);

    input E;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $_OAI4_
(
    D,
    C,
    B,
    A,
    Y
);

    input D;
    input C;
    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $_AOI4_
(
    D,
    C,
    B,
    A,
    Y
);

    input D;
    input C;
    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $_OAI3_
(
    C,
    B,
    A,
    Y
);

    input C;
    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $_AOI3_
(
    C,
    B,
    A,
    Y
);

    input C;
    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $_MUX16_
(
    V,
    U,
    T,
    S,
    P,
    O,
    N,
    M,
    L,
    K,
    J,
    I,
    H,
    G,
    F,
    E,
    D,
    C,
    B,
    A,
    Y
);

    input V;
    input U;
    input T;
    input S;
    input P;
    input O;
    input N;
    input M;
    input L;
    input K;
    input J;
    input I;
    input H;
    input G;
    input F;
    input E;
    input D;
    input C;
    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $_MUX8_
(
    U,
    T,
    S,
    H,
    G,
    F,
    E,
    D,
    C,
    B,
    A,
    Y
);

    input U;
    input T;
    input S;
    input H;
    input G;
    input F;
    input E;
    input D;
    input C;
    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $_MUX4_
(
    T,
    S,
    D,
    C,
    B,
    A,
    Y
);

    input T;
    input S;
    input D;
    input C;
    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $_NMUX_
(
    S,
    B,
    A,
    Y
);

    input S;
    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $_MUX_
(
    S,
    B,
    A,
    Y
);

    input S;
    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $_ORNOT_
(
    B,
    A,
    Y
);

    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $_ANDNOT_
(
    B,
    A,
    Y
);

    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $_XNOR_
(
    B,
    A,
    Y
);

    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $_XOR_
(
    B,
    A,
    Y
);

    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $_NOR_
(
    B,
    A,
    Y
);

    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $_OR_
(
    B,
    A,
    Y
);

    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $_NAND_
(
    B,
    A,
    Y
);

    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $_AND_
(
    B,
    A,
    Y
);

    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $_NOT_
(
    A,
    Y
);

    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $_BUF_
(
    A,
    Y
);

    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $fsm
(
    CTRL_IN,
    ARST,
    CLK,
    CTRL_OUT
);

    input CTRL_IN;
    input ARST;
    input CLK;
    output CTRL_OUT;

endmodule
`endcelldefine

`celldefine
module $mem_v2
(
    WR_DATA,
    WR_ADDR,
    WR_EN,
    WR_CLK,
    RD_ADDR,
    RD_SRST,
    RD_ARST,
    RD_EN,
    RD_CLK,
    RD_DATA
);

    input WR_DATA;
    input WR_ADDR;
    input WR_EN;
    input WR_CLK;
    input RD_ADDR;
    input RD_SRST;
    input RD_ARST;
    input RD_EN;
    input RD_CLK;
    output RD_DATA;

endmodule
`endcelldefine

`celldefine
module $mem
(
    WR_DATA,
    WR_ADDR,
    WR_EN,
    WR_CLK,
    RD_ADDR,
    RD_EN,
    RD_CLK,
    RD_DATA
);

    input WR_DATA;
    input WR_ADDR;
    input WR_EN;
    input WR_CLK;
    input RD_ADDR;
    input RD_EN;
    input RD_CLK;
    output RD_DATA;

endmodule
`endcelldefine

`celldefine
module $meminit_v2
(
    EN,
    DATA,
    ADDR
);

    input EN;
    input DATA;
    input ADDR;

endmodule
`endcelldefine

`celldefine
module $meminit
(
    DATA,
    ADDR
);

    input DATA;
    input ADDR;

endmodule
`endcelldefine

`celldefine
module $memwr_v2
(
    DATA,
    ADDR,
    EN,
    CLK
);

    input DATA;
    input ADDR;
    input EN;
    input CLK;

endmodule
`endcelldefine

`celldefine
module $memwr
(
    DATA,
    ADDR,
    EN,
    CLK
);

    input DATA;
    input ADDR;
    input EN;
    input CLK;

endmodule
`endcelldefine

`celldefine
module $memrd_v2
(
    ADDR,
    SRST,
    ARST,
    EN,
    CLK,
    DATA
);

    input ADDR;
    input SRST;
    input ARST;
    input EN;
    input CLK;
    output DATA;

endmodule
`endcelldefine

`celldefine
module $memrd
(
    ADDR,
    EN,
    CLK,
    DATA
);

    input ADDR;
    input EN;
    input CLK;
    output DATA;

endmodule
`endcelldefine

`celldefine
module $dlatchsr
(
    D,
    CLR,
    SET,
    EN,
    Q
);

    input D;
    input CLR;
    input SET;
    input EN;
    output Q;

endmodule
`endcelldefine

`celldefine
module $adlatch
(
    ARST,
    D,
    EN,
    Q
);

    input ARST;
    input D;
    input EN;
    output Q;

endmodule
`endcelldefine

`celldefine
module $dlatch
(
    D,
    EN,
    Q
);

    input D;
    input EN;
    output Q;

endmodule
`endcelldefine

`celldefine
module $sdffce
(
    EN,
    D,
    SRST,
    CLK,
    Q
);

    input EN;
    input D;
    input SRST;
    input CLK;
    output Q;

endmodule
`endcelldefine

`celldefine
module $sdffe
(
    EN,
    D,
    SRST,
    CLK,
    Q
);

    input EN;
    input D;
    input SRST;
    input CLK;
    output Q;

endmodule
`endcelldefine

`celldefine
module $sdff
(
    D,
    SRST,
    CLK,
    Q
);

    input D;
    input SRST;
    input CLK;
    output Q;

endmodule
`endcelldefine

`celldefine
module $aldffe
(
    EN,
    D,
    AD,
    ALOAD,
    CLK,
    Q
);

    input EN;
    input D;
    input AD;
    input ALOAD;
    input CLK;
    output Q;

endmodule
`endcelldefine

`celldefine
module $aldff
(
    D,
    AD,
    ALOAD,
    CLK,
    Q
);

    input D;
    input AD;
    input ALOAD;
    input CLK;
    output Q;

endmodule
`endcelldefine

`celldefine
module $adffe
(
    EN,
    D,
    ARST,
    CLK,
    Q
);

    input EN;
    input D;
    input ARST;
    input CLK;
    output Q;

endmodule
`endcelldefine

`celldefine
module $adff
(
    D,
    ARST,
    CLK,
    Q
);

    input D;
    input ARST;
    input CLK;
    output Q;

endmodule
`endcelldefine

`celldefine
module $dffsre
(
    EN,
    D,
    CLR,
    SET,
    CLK,
    Q
);

    input EN;
    input D;
    input CLR;
    input SET;
    input CLK;
    output Q;

endmodule
`endcelldefine

`celldefine
module $dffsr
(
    D,
    CLR,
    SET,
    CLK,
    Q
);

    input D;
    input CLR;
    input SET;
    input CLK;
    output Q;

endmodule
`endcelldefine

`celldefine
module $dffe
(
    D,
    EN,
    CLK,
    Q
);

    input D;
    input EN;
    input CLK;
    output Q;

endmodule
`endcelldefine

`celldefine
module $dff
(
    D,
    CLK,
    Q
);

    input D;
    input CLK;
    output Q;

endmodule
`endcelldefine

`celldefine
module $ff
(
    D,
    Q
);

    input D;
    output Q;

endmodule
`endcelldefine

`celldefine
module $sr
(
    CLR,
    SET,
    Q
);

    input CLR;
    input SET;
    output Q;

endmodule
`endcelldefine

`celldefine
module $specrule
(
    DST,
    SRC,
    EN_DST,
    EN_SRC
);

    input DST;
    input SRC;
    input EN_DST;
    input EN_SRC;

endmodule
`endcelldefine

`celldefine
module $specify3
(
    DAT,
    DST,
    SRC,
    EN
);

    input DAT;
    input DST;
    input SRC;
    input EN;

endmodule
`endcelldefine

`celldefine
module $specify2
(
    DST,
    SRC,
    EN
);

    input DST;
    input SRC;
    input EN;

endmodule
`endcelldefine

`celldefine
module $equiv
(
    B,
    A,
    Y
);

    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $allseq
(
    Y
);

    output Y;

endmodule
`endcelldefine

`celldefine
module $allconst
(
    Y
);

    output Y;

endmodule
`endcelldefine

`celldefine
module $anyseq
(
    Y
);

    output Y;

endmodule
`endcelldefine

`celldefine
module $anyconst
(
    Y
);

    output Y;

endmodule
`endcelldefine

`celldefine
module $initstate
(
    Y
);

    output Y;

endmodule
`endcelldefine

`celldefine
module $cover
(
    EN,
    A
);

    input EN;
    input A;

endmodule
`endcelldefine

`celldefine
module $fair
(
    EN,
    A
);

    input EN;
    input A;

endmodule
`endcelldefine

`celldefine
module $live
(
    EN,
    A
);

    input EN;
    input A;

endmodule
`endcelldefine

`celldefine
module $assume
(
    EN,
    A
);

    input EN;
    input A;

endmodule
`endcelldefine

`celldefine
module $assert
(
    EN,
    A
);

    input EN;
    input A;

endmodule
`endcelldefine

`celldefine
module $tribuf
(
    EN,
    A,
    Y
);

    input EN;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $fa
(
    C,
    B,
    A,
    Y,
    X
);

    input C;
    input B;
    input A;
    output Y;
    output X;

endmodule
`endcelldefine

`celldefine
module $alu
(
    BI,
    CI,
    B,
    A,
    CO,
    Y,
    X
);

    input BI;
    input CI;
    input B;
    input A;
    output CO;
    output Y;
    output X;

endmodule
`endcelldefine

`celldefine
module $lcu
(
    CI,
    G,
    P,
    CO
);

    input CI;
    input G;
    input P;
    output CO;

endmodule
`endcelldefine

`celldefine
module $demux
(
    S,
    A,
    Y
);

    input S;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $bmux
(
    S,
    A,
    Y
);

    input S;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $pmux
(
    S,
    B,
    A,
    Y
);

    input S;
    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $mux
(
    S,
    B,
    A,
    Y
);

    input S;
    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $macc
(
    B,
    A,
    Y
);

    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $concat
(
    B,
    A,
    Y
);

    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $logic_or
(
    B,
    A,
    Y
);

    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $logic_and
(
    B,
    A,
    Y
);

    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $pow
(
    B,
    A,
    Y
);

    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $modfloor
(
    B,
    A,
    Y
);

    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $divfloor
(
    B,
    A,
    Y
);

    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $mod
(
    B,
    A,
    Y
);

    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $div
(
    B,
    A,
    Y
);

    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $mul
(
    B,
    A,
    Y
);

    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $sub
(
    B,
    A,
    Y
);

    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $add
(
    B,
    A,
    Y
);

    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $gt
(
    B,
    A,
    Y
);

    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $ge
(
    B,
    A,
    Y
);

    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $nex
(
    B,
    A,
    Y
);

    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $eqx
(
    B,
    A,
    Y
);

    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $ne
(
    B,
    A,
    Y
);

    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $eq
(
    B,
    A,
    Y
);

    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $le
(
    B,
    A,
    Y
);

    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $lt
(
    B,
    A,
    Y
);

    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $shiftx
(
    B,
    A,
    Y
);

    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $shift
(
    B,
    A,
    Y
);

    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $sshr
(
    B,
    A,
    Y
);

    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $sshl
(
    B,
    A,
    Y
);

    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $shr
(
    B,
    A,
    Y
);

    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $shl
(
    B,
    A,
    Y
);

    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $xnor
(
    B,
    A,
    Y
);

    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $xor
(
    B,
    A,
    Y
);

    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $or
(
    B,
    A,
    Y
);

    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $and
(
    B,
    A,
    Y
);

    input B;
    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $sop
(
    A,
    Y
);

    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $lut
(
    A,
    Y
);

    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $slice
(
    A,
    Y
);

    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $logic_not
(
    A,
    Y
);

    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $reduce_bool
(
    A,
    Y
);

    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $reduce_xnor
(
    A,
    Y
);

    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $reduce_xor
(
    A,
    Y
);

    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $reduce_or
(
    A,
    Y
);

    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $reduce_and
(
    A,
    Y
);

    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $neg
(
    A,
    Y
);

    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $pos
(
    A,
    Y
);

    input A;
    output Y;

endmodule
`endcelldefine

`celldefine
module $not
(
    A,
    Y
);

    input A;
    output Y;

endmodule
`endcelldefine

