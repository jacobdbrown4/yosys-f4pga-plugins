module not_ft(
    A_TMR_0,
    A_TMR_1,
    A_TMR_2,
    Y_TMR_0,
    Y_TMR_1,
    Y_TMR_2
);

    parameter A_SIGNED = 0;
    parameter A_WIDTH  = 1;
    parameter Y_WIDTH = 1;

    input A_TMR_0;
    input A_TMR_1;
    input A_TMR_2;
    output Y_TMR_0;
    output Y_TMR_1;
    output Y_TMR_2;

endmodule